module main_0
   (IN1_STB,
    OUT1_ACK,
    E,
    DATA_ACK,
    Q,
    ETH_CLK_OBUF,
    INTERNAL_RST_reg,
    S_IN1_ACK_reg,
    OUT1_STB_reg,
    S_DATA_STB_reg,
    OUT1_STB,
    DATA,
    OUT1,
    IN1_ACK,
    S_DATA_STB_reg_0);
  output IN1_STB;
  output OUT1_ACK;
  output [0:0]E;
  output DATA_ACK;
  output [7:0]Q;
  input ETH_CLK_OBUF;
  input INTERNAL_RST_reg;
  input S_IN1_ACK_reg;
  input OUT1_STB_reg;
  input S_DATA_STB_reg;
  input OUT1_STB;
  input [7:0]DATA;
  input [7:0]OUT1;
  input IN1_ACK;
  input S_DATA_STB_reg_0;
  wire [7:0]DATA;
  wire DATA_ACK;
  wire [0:0]E;
  wire ETH_CLK_OBUF;
  wire IN1_ACK;
  wire IN1_STB;
  wire INTERNAL_RST_reg;
  wire [7:0]OUT1;
  wire OUT1_ACK;
  wire OUT1_STB;
  wire OUT1_STB_reg;
  wire [7:0]Q;
  wire S_DATA_STB_reg;
  wire S_DATA_STB_reg_0;
  wire S_IN1_ACK_reg;
  wire [3:0]address_a;
  wire [3:0]address_a_2;
  wire [3:0]address_b_2;
  wire [3:0]address_z;
  wire [3:0]address_z_2;
  wire [3:0]address_z_3;
  wire \address_z_3[3]_i_1_n_0 ;
  wire [15:1]data1;
  wire [16:1]data2;
  wire [31:0]data4;
  wire [31:0]data5;
  wire instruction0;
  wire \instruction[0]_i_11_n_0 ;
  wire \instruction[0]_i_12_n_0 ;
  wire \instruction[0]_i_13_n_0 ;
  wire \instruction[0]_i_14_n_0 ;
  wire \instruction[0]_i_15_n_0 ;
  wire \instruction[0]_i_16_n_0 ;
  wire \instruction[0]_i_17_n_0 ;
  wire \instruction[0]_i_18_n_0 ;
  wire \instruction[0]_i_19_n_0 ;
  wire \instruction[0]_i_1_n_0 ;
  wire \instruction[0]_i_21_n_0 ;
  wire \instruction[0]_i_22_n_0 ;
  wire \instruction[0]_i_23_n_0 ;
  wire \instruction[0]_i_25_n_0 ;
  wire \instruction[0]_i_26_n_0 ;
  wire \instruction[0]_i_28_n_0 ;
  wire \instruction[0]_i_29_n_0 ;
  wire \instruction[0]_i_30_n_0 ;
  wire \instruction[0]_i_31_n_0 ;
  wire \instruction[0]_i_32_n_0 ;
  wire \instruction[0]_i_34_n_0 ;
  wire \instruction[0]_i_35_n_0 ;
  wire \instruction[0]_i_38_n_0 ;
  wire \instruction[0]_i_3_n_0 ;
  wire \instruction[0]_i_40_n_0 ;
  wire \instruction[0]_i_41_n_0 ;
  wire \instruction[0]_i_42_n_0 ;
  wire \instruction[0]_i_43_n_0 ;
  wire \instruction[0]_i_44_n_0 ;
  wire \instruction[0]_i_45_n_0 ;
  wire \instruction[0]_i_46_n_0 ;
  wire \instruction[0]_i_48_n_0 ;
  wire \instruction[0]_i_49_n_0 ;
  wire \instruction[0]_i_51_n_0 ;
  wire \instruction[0]_i_52_n_0 ;
  wire \instruction[0]_i_53_n_0 ;
  wire \instruction[0]_i_54_n_0 ;
  wire \instruction[0]_i_55_n_0 ;
  wire \instruction[0]_i_56_n_0 ;
  wire \instruction[0]_i_57_n_0 ;
  wire \instruction[0]_i_58_n_0 ;
  wire \instruction[0]_i_59_n_0 ;
  wire \instruction[0]_i_60_n_0 ;
  wire \instruction[0]_i_61_n_0 ;
  wire \instruction[0]_i_62_n_0 ;
  wire \instruction[0]_i_63_n_0 ;
  wire \instruction[0]_i_6_n_0 ;
  wire \instruction[0]_i_7_n_0 ;
  wire \instruction[0]_i_8_n_0 ;
  wire \instruction[0]_i_9_n_0 ;
  wire \instruction[15]_i_10_n_0 ;
  wire \instruction[15]_i_11_n_0 ;
  wire \instruction[15]_i_12_n_0 ;
  wire \instruction[15]_i_13_n_0 ;
  wire \instruction[15]_i_14_n_0 ;
  wire \instruction[15]_i_15_n_0 ;
  wire \instruction[15]_i_16_n_0 ;
  wire \instruction[15]_i_17_n_0 ;
  wire \instruction[15]_i_18_n_0 ;
  wire \instruction[15]_i_1_n_0 ;
  wire \instruction[15]_i_2_n_0 ;
  wire \instruction[15]_i_3_n_0 ;
  wire \instruction[15]_i_4_n_0 ;
  wire \instruction[15]_i_5_n_0 ;
  wire \instruction[15]_i_6_n_0 ;
  wire \instruction[15]_i_7_n_0 ;
  wire \instruction[15]_i_8_n_0 ;
  wire \instruction[15]_i_9_n_0 ;
  wire \instruction[16]_i_10_n_0 ;
  wire \instruction[16]_i_11_n_0 ;
  wire \instruction[16]_i_12_n_0 ;
  wire \instruction[16]_i_13_n_0 ;
  wire \instruction[16]_i_14_n_0 ;
  wire \instruction[16]_i_15_n_0 ;
  wire \instruction[16]_i_16_n_0 ;
  wire \instruction[16]_i_19_n_0 ;
  wire \instruction[16]_i_1_n_0 ;
  wire \instruction[16]_i_20_n_0 ;
  wire \instruction[16]_i_21_n_0 ;
  wire \instruction[16]_i_23_n_0 ;
  wire \instruction[16]_i_24_n_0 ;
  wire \instruction[16]_i_25_n_0 ;
  wire \instruction[16]_i_26_n_0 ;
  wire \instruction[16]_i_27_n_0 ;
  wire \instruction[16]_i_28_n_0 ;
  wire \instruction[16]_i_29_n_0 ;
  wire \instruction[16]_i_2_n_0 ;
  wire \instruction[16]_i_30_n_0 ;
  wire \instruction[16]_i_31_n_0 ;
  wire \instruction[16]_i_32_n_0 ;
  wire \instruction[16]_i_33_n_0 ;
  wire \instruction[16]_i_34_n_0 ;
  wire \instruction[16]_i_35_n_0 ;
  wire \instruction[16]_i_36_n_0 ;
  wire \instruction[16]_i_37_n_0 ;
  wire \instruction[16]_i_38_n_0 ;
  wire \instruction[16]_i_39_n_0 ;
  wire \instruction[16]_i_40_n_0 ;
  wire \instruction[16]_i_41_n_0 ;
  wire \instruction[16]_i_42_n_0 ;
  wire \instruction[16]_i_43_n_0 ;
  wire \instruction[16]_i_44_n_0 ;
  wire \instruction[16]_i_45_n_0 ;
  wire \instruction[16]_i_4_n_0 ;
  wire \instruction[16]_i_6_n_0 ;
  wire \instruction[16]_i_7_n_0 ;
  wire \instruction[16]_i_8_n_0 ;
  wire \instruction[16]_i_9_n_0 ;
  wire \instruction[17]_i_10_n_0 ;
  wire \instruction[17]_i_11_n_0 ;
  wire \instruction[17]_i_13_n_0 ;
  wire \instruction[17]_i_15_n_0 ;
  wire \instruction[17]_i_16_n_0 ;
  wire \instruction[17]_i_17_n_0 ;
  wire \instruction[17]_i_18_n_0 ;
  wire \instruction[17]_i_19_n_0 ;
  wire \instruction[17]_i_1_n_0 ;
  wire \instruction[17]_i_20_n_0 ;
  wire \instruction[17]_i_21_n_0 ;
  wire \instruction[17]_i_22_n_0 ;
  wire \instruction[17]_i_23_n_0 ;
  wire \instruction[17]_i_24_n_0 ;
  wire \instruction[17]_i_25_n_0 ;
  wire \instruction[17]_i_27_n_0 ;
  wire \instruction[17]_i_28_n_0 ;
  wire \instruction[17]_i_29_n_0 ;
  wire \instruction[17]_i_2_n_0 ;
  wire \instruction[17]_i_31_n_0 ;
  wire \instruction[17]_i_32_n_0 ;
  wire \instruction[17]_i_33_n_0 ;
  wire \instruction[17]_i_34_n_0 ;
  wire \instruction[17]_i_35_n_0 ;
  wire \instruction[17]_i_36_n_0 ;
  wire \instruction[17]_i_37_n_0 ;
  wire \instruction[17]_i_38_n_0 ;
  wire \instruction[17]_i_39_n_0 ;
  wire \instruction[17]_i_40_n_0 ;
  wire \instruction[17]_i_41_n_0 ;
  wire \instruction[17]_i_42_n_0 ;
  wire \instruction[17]_i_43_n_0 ;
  wire \instruction[17]_i_44_n_0 ;
  wire \instruction[17]_i_45_n_0 ;
  wire \instruction[17]_i_47_n_0 ;
  wire \instruction[17]_i_48_n_0 ;
  wire \instruction[17]_i_49_n_0 ;
  wire \instruction[17]_i_50_n_0 ;
  wire \instruction[17]_i_51_n_0 ;
  wire \instruction[17]_i_5_n_0 ;
  wire \instruction[17]_i_6_n_0 ;
  wire \instruction[17]_i_7_n_0 ;
  wire \instruction[17]_i_8_n_0 ;
  wire \instruction[17]_i_9_n_0 ;
  wire \instruction[18]_i_11_n_0 ;
  wire \instruction[18]_i_14_n_0 ;
  wire \instruction[18]_i_15_n_0 ;
  wire \instruction[18]_i_16_n_0 ;
  wire \instruction[18]_i_17_n_0 ;
  wire \instruction[18]_i_18_n_0 ;
  wire \instruction[18]_i_19_n_0 ;
  wire \instruction[18]_i_1_n_0 ;
  wire \instruction[18]_i_20_n_0 ;
  wire \instruction[18]_i_24_n_0 ;
  wire \instruction[18]_i_25_n_0 ;
  wire \instruction[18]_i_26_n_0 ;
  wire \instruction[18]_i_27_n_0 ;
  wire \instruction[18]_i_28_n_0 ;
  wire \instruction[18]_i_29_n_0 ;
  wire \instruction[18]_i_2_n_0 ;
  wire \instruction[18]_i_30_n_0 ;
  wire \instruction[18]_i_31_n_0 ;
  wire \instruction[18]_i_32_n_0 ;
  wire \instruction[18]_i_33_n_0 ;
  wire \instruction[18]_i_34_n_0 ;
  wire \instruction[18]_i_35_n_0 ;
  wire \instruction[18]_i_36_n_0 ;
  wire \instruction[18]_i_37_n_0 ;
  wire \instruction[18]_i_38_n_0 ;
  wire \instruction[18]_i_39_n_0 ;
  wire \instruction[18]_i_3_n_0 ;
  wire \instruction[18]_i_40_n_0 ;
  wire \instruction[18]_i_41_n_0 ;
  wire \instruction[18]_i_42_n_0 ;
  wire \instruction[18]_i_6_n_0 ;
  wire \instruction[18]_i_7_n_0 ;
  wire \instruction[18]_i_9_n_0 ;
  wire \instruction[19]_i_11_n_0 ;
  wire \instruction[19]_i_13_n_0 ;
  wire \instruction[19]_i_14_n_0 ;
  wire \instruction[19]_i_15_n_0 ;
  wire \instruction[19]_i_16_n_0 ;
  wire \instruction[19]_i_17_n_0 ;
  wire \instruction[19]_i_18_n_0 ;
  wire \instruction[19]_i_19_n_0 ;
  wire \instruction[19]_i_1_n_0 ;
  wire \instruction[19]_i_20_n_0 ;
  wire \instruction[19]_i_21_n_0 ;
  wire \instruction[19]_i_22_n_0 ;
  wire \instruction[19]_i_23_n_0 ;
  wire \instruction[19]_i_24_n_0 ;
  wire \instruction[19]_i_25_n_0 ;
  wire \instruction[19]_i_26_n_0 ;
  wire \instruction[19]_i_27_n_0 ;
  wire \instruction[19]_i_28_n_0 ;
  wire \instruction[19]_i_29_n_0 ;
  wire \instruction[19]_i_2_n_0 ;
  wire \instruction[19]_i_30_n_0 ;
  wire \instruction[19]_i_31_n_0 ;
  wire \instruction[19]_i_32_n_0 ;
  wire \instruction[19]_i_3_n_0 ;
  wire \instruction[19]_i_4_n_0 ;
  wire \instruction[19]_i_5_n_0 ;
  wire \instruction[19]_i_6_n_0 ;
  wire \instruction[19]_i_7_n_0 ;
  wire \instruction[19]_i_8_n_0 ;
  wire \instruction[19]_i_9_n_0 ;
  wire \instruction[1]_i_10_n_0 ;
  wire \instruction[1]_i_11_n_0 ;
  wire \instruction[1]_i_12_n_0 ;
  wire \instruction[1]_i_13_n_0 ;
  wire \instruction[1]_i_14_n_0 ;
  wire \instruction[1]_i_15_n_0 ;
  wire \instruction[1]_i_16_n_0 ;
  wire \instruction[1]_i_19_n_0 ;
  wire \instruction[1]_i_1_n_0 ;
  wire \instruction[1]_i_20_n_0 ;
  wire \instruction[1]_i_21_n_0 ;
  wire \instruction[1]_i_22_n_0 ;
  wire \instruction[1]_i_25_n_0 ;
  wire \instruction[1]_i_26_n_0 ;
  wire \instruction[1]_i_27_n_0 ;
  wire \instruction[1]_i_28_n_0 ;
  wire \instruction[1]_i_29_n_0 ;
  wire \instruction[1]_i_30_n_0 ;
  wire \instruction[1]_i_31_n_0 ;
  wire \instruction[1]_i_32_n_0 ;
  wire \instruction[1]_i_33_n_0 ;
  wire \instruction[1]_i_34_n_0 ;
  wire \instruction[1]_i_35_n_0 ;
  wire \instruction[1]_i_36_n_0 ;
  wire \instruction[1]_i_37_n_0 ;
  wire \instruction[1]_i_38_n_0 ;
  wire \instruction[1]_i_39_n_0 ;
  wire \instruction[1]_i_3_n_0 ;
  wire \instruction[1]_i_40_n_0 ;
  wire \instruction[1]_i_41_n_0 ;
  wire \instruction[1]_i_42_n_0 ;
  wire \instruction[1]_i_43_n_0 ;
  wire \instruction[1]_i_44_n_0 ;
  wire \instruction[1]_i_45_n_0 ;
  wire \instruction[1]_i_46_n_0 ;
  wire \instruction[1]_i_47_n_0 ;
  wire \instruction[1]_i_49_n_0 ;
  wire \instruction[1]_i_51_n_0 ;
  wire \instruction[1]_i_54_n_0 ;
  wire \instruction[1]_i_55_n_0 ;
  wire \instruction[1]_i_56_n_0 ;
  wire \instruction[1]_i_57_n_0 ;
  wire \instruction[1]_i_58_n_0 ;
  wire \instruction[1]_i_59_n_0 ;
  wire \instruction[1]_i_60_n_0 ;
  wire \instruction[1]_i_61_n_0 ;
  wire \instruction[1]_i_8_n_0 ;
  wire \instruction[1]_i_9_n_0 ;
  wire \instruction[20]_i_10_n_0 ;
  wire \instruction[20]_i_11_n_0 ;
  wire \instruction[20]_i_13_n_0 ;
  wire \instruction[20]_i_14_n_0 ;
  wire \instruction[20]_i_15_n_0 ;
  wire \instruction[20]_i_16_n_0 ;
  wire \instruction[20]_i_17_n_0 ;
  wire \instruction[20]_i_18_n_0 ;
  wire \instruction[20]_i_19_n_0 ;
  wire \instruction[20]_i_1_n_0 ;
  wire \instruction[20]_i_20_n_0 ;
  wire \instruction[20]_i_21_n_0 ;
  wire \instruction[20]_i_22_n_0 ;
  wire \instruction[20]_i_24_n_0 ;
  wire \instruction[20]_i_26_n_0 ;
  wire \instruction[20]_i_27_n_0 ;
  wire \instruction[20]_i_28_n_0 ;
  wire \instruction[20]_i_29_n_0 ;
  wire \instruction[20]_i_2_n_0 ;
  wire \instruction[20]_i_30_n_0 ;
  wire \instruction[20]_i_31_n_0 ;
  wire \instruction[20]_i_3_n_0 ;
  wire \instruction[20]_i_4_n_0 ;
  wire \instruction[20]_i_5_n_0 ;
  wire \instruction[20]_i_6_n_0 ;
  wire \instruction[20]_i_7_n_0 ;
  wire \instruction[20]_i_9_n_0 ;
  wire \instruction[21]_i_12_n_0 ;
  wire \instruction[21]_i_14_n_0 ;
  wire \instruction[21]_i_15_n_0 ;
  wire \instruction[21]_i_16_n_0 ;
  wire \instruction[21]_i_17_n_0 ;
  wire \instruction[21]_i_18_n_0 ;
  wire \instruction[21]_i_19_n_0 ;
  wire \instruction[21]_i_1_n_0 ;
  wire \instruction[21]_i_20_n_0 ;
  wire \instruction[21]_i_21_n_0 ;
  wire \instruction[21]_i_22_n_0 ;
  wire \instruction[21]_i_23_n_0 ;
  wire \instruction[21]_i_24_n_0 ;
  wire \instruction[21]_i_25_n_0 ;
  wire \instruction[21]_i_26_n_0 ;
  wire \instruction[21]_i_27_n_0 ;
  wire \instruction[21]_i_28_n_0 ;
  wire \instruction[21]_i_29_n_0 ;
  wire \instruction[21]_i_2_n_0 ;
  wire \instruction[21]_i_30_n_0 ;
  wire \instruction[21]_i_31_n_0 ;
  wire \instruction[21]_i_32_n_0 ;
  wire \instruction[21]_i_37_n_0 ;
  wire \instruction[21]_i_38_n_0 ;
  wire \instruction[21]_i_3_n_0 ;
  wire \instruction[21]_i_41_n_0 ;
  wire \instruction[21]_i_42_n_0 ;
  wire \instruction[21]_i_43_n_0 ;
  wire \instruction[21]_i_45_n_0 ;
  wire \instruction[21]_i_46_n_0 ;
  wire \instruction[21]_i_47_n_0 ;
  wire \instruction[21]_i_48_n_0 ;
  wire \instruction[21]_i_49_n_0 ;
  wire \instruction[21]_i_50_n_0 ;
  wire \instruction[21]_i_51_n_0 ;
  wire \instruction[21]_i_52_n_0 ;
  wire \instruction[21]_i_53_n_0 ;
  wire \instruction[21]_i_54_n_0 ;
  wire \instruction[21]_i_55_n_0 ;
  wire \instruction[21]_i_56_n_0 ;
  wire \instruction[21]_i_57_n_0 ;
  wire \instruction[21]_i_58_n_0 ;
  wire \instruction[21]_i_59_n_0 ;
  wire \instruction[21]_i_60_n_0 ;
  wire \instruction[21]_i_61_n_0 ;
  wire \instruction[21]_i_62_n_0 ;
  wire \instruction[21]_i_63_n_0 ;
  wire \instruction[21]_i_6_n_0 ;
  wire \instruction[21]_i_7_n_0 ;
  wire \instruction[21]_i_8_n_0 ;
  wire \instruction[21]_i_9_n_0 ;
  wire \instruction[22]_i_10_n_0 ;
  wire \instruction[22]_i_11_n_0 ;
  wire \instruction[22]_i_12_n_0 ;
  wire \instruction[22]_i_13_n_0 ;
  wire \instruction[22]_i_1_n_0 ;
  wire \instruction[22]_i_2_n_0 ;
  wire \instruction[22]_i_3_n_0 ;
  wire \instruction[22]_i_4_n_0 ;
  wire \instruction[22]_i_6_n_0 ;
  wire \instruction[22]_i_7_n_0 ;
  wire \instruction[22]_i_8_n_0 ;
  wire \instruction[22]_i_9_n_0 ;
  wire \instruction[23]_i_11_n_0 ;
  wire \instruction[23]_i_12_n_0 ;
  wire \instruction[23]_i_13_n_0 ;
  wire \instruction[23]_i_14_n_0 ;
  wire \instruction[23]_i_15_n_0 ;
  wire \instruction[23]_i_16_n_0 ;
  wire \instruction[23]_i_17_n_0 ;
  wire \instruction[23]_i_18_n_0 ;
  wire \instruction[23]_i_19_n_0 ;
  wire \instruction[23]_i_1_n_0 ;
  wire \instruction[23]_i_20_n_0 ;
  wire \instruction[23]_i_21_n_0 ;
  wire \instruction[23]_i_22_n_0 ;
  wire \instruction[23]_i_23_n_0 ;
  wire \instruction[23]_i_24_n_0 ;
  wire \instruction[23]_i_25_n_0 ;
  wire \instruction[23]_i_26_n_0 ;
  wire \instruction[23]_i_28_n_0 ;
  wire \instruction[23]_i_29_n_0 ;
  wire \instruction[23]_i_30_n_0 ;
  wire \instruction[23]_i_31_n_0 ;
  wire \instruction[23]_i_32_n_0 ;
  wire \instruction[23]_i_34_n_0 ;
  wire \instruction[23]_i_35_n_0 ;
  wire \instruction[23]_i_36_n_0 ;
  wire \instruction[23]_i_37_n_0 ;
  wire \instruction[23]_i_38_n_0 ;
  wire \instruction[23]_i_39_n_0 ;
  wire \instruction[23]_i_3_n_0 ;
  wire \instruction[23]_i_41_n_0 ;
  wire \instruction[23]_i_42_n_0 ;
  wire \instruction[23]_i_46_n_0 ;
  wire \instruction[23]_i_47_n_0 ;
  wire \instruction[23]_i_48_n_0 ;
  wire \instruction[23]_i_49_n_0 ;
  wire \instruction[23]_i_50_n_0 ;
  wire \instruction[23]_i_51_n_0 ;
  wire \instruction[23]_i_52_n_0 ;
  wire \instruction[23]_i_53_n_0 ;
  wire \instruction[23]_i_54_n_0 ;
  wire \instruction[23]_i_55_n_0 ;
  wire \instruction[23]_i_56_n_0 ;
  wire \instruction[23]_i_57_n_0 ;
  wire \instruction[23]_i_7_n_0 ;
  wire \instruction[23]_i_8_n_0 ;
  wire \instruction[23]_i_9_n_0 ;
  wire \instruction[24]_i_10_n_0 ;
  wire \instruction[24]_i_11_n_0 ;
  wire \instruction[24]_i_12_n_0 ;
  wire \instruction[24]_i_13_n_0 ;
  wire \instruction[24]_i_14_n_0 ;
  wire \instruction[24]_i_15_n_0 ;
  wire \instruction[24]_i_16_n_0 ;
  wire \instruction[24]_i_17_n_0 ;
  wire \instruction[24]_i_18_n_0 ;
  wire \instruction[24]_i_1_n_0 ;
  wire \instruction[24]_i_21_n_0 ;
  wire \instruction[24]_i_22_n_0 ;
  wire \instruction[24]_i_23_n_0 ;
  wire \instruction[24]_i_24_n_0 ;
  wire \instruction[24]_i_26_n_0 ;
  wire \instruction[24]_i_27_n_0 ;
  wire \instruction[24]_i_28_n_0 ;
  wire \instruction[24]_i_29_n_0 ;
  wire \instruction[24]_i_2_n_0 ;
  wire \instruction[24]_i_30_n_0 ;
  wire \instruction[24]_i_31_n_0 ;
  wire \instruction[24]_i_32_n_0 ;
  wire \instruction[24]_i_33_n_0 ;
  wire \instruction[24]_i_34_n_0 ;
  wire \instruction[24]_i_35_n_0 ;
  wire \instruction[24]_i_36_n_0 ;
  wire \instruction[24]_i_37_n_0 ;
  wire \instruction[24]_i_38_n_0 ;
  wire \instruction[24]_i_39_n_0 ;
  wire \instruction[24]_i_40_n_0 ;
  wire \instruction[24]_i_42_n_0 ;
  wire \instruction[24]_i_43_n_0 ;
  wire \instruction[24]_i_44_n_0 ;
  wire \instruction[24]_i_46_n_0 ;
  wire \instruction[24]_i_47_n_0 ;
  wire \instruction[24]_i_48_n_0 ;
  wire \instruction[24]_i_49_n_0 ;
  wire \instruction[24]_i_50_n_0 ;
  wire \instruction[24]_i_51_n_0 ;
  wire \instruction[24]_i_52_n_0 ;
  wire \instruction[24]_i_53_n_0 ;
  wire \instruction[24]_i_54_n_0 ;
  wire \instruction[24]_i_55_n_0 ;
  wire \instruction[24]_i_56_n_0 ;
  wire \instruction[24]_i_57_n_0 ;
  wire \instruction[24]_i_6_n_0 ;
  wire \instruction[24]_i_7_n_0 ;
  wire \instruction[24]_i_8_n_0 ;
  wire \instruction[24]_i_9_n_0 ;
  wire \instruction[25]_i_10_n_0 ;
  wire \instruction[25]_i_11_n_0 ;
  wire \instruction[25]_i_12_n_0 ;
  wire \instruction[25]_i_13_n_0 ;
  wire \instruction[25]_i_14_n_0 ;
  wire \instruction[25]_i_15_n_0 ;
  wire \instruction[25]_i_16_n_0 ;
  wire \instruction[25]_i_17_n_0 ;
  wire \instruction[25]_i_18_n_0 ;
  wire \instruction[25]_i_1_n_0 ;
  wire \instruction[25]_i_21_n_0 ;
  wire \instruction[25]_i_22_n_0 ;
  wire \instruction[25]_i_23_n_0 ;
  wire \instruction[25]_i_24_n_0 ;
  wire \instruction[25]_i_25_n_0 ;
  wire \instruction[25]_i_27_n_0 ;
  wire \instruction[25]_i_28_n_0 ;
  wire \instruction[25]_i_29_n_0 ;
  wire \instruction[25]_i_2_n_0 ;
  wire \instruction[25]_i_30_n_0 ;
  wire \instruction[25]_i_35_n_0 ;
  wire \instruction[25]_i_36_n_0 ;
  wire \instruction[25]_i_37_n_0 ;
  wire \instruction[25]_i_38_n_0 ;
  wire \instruction[25]_i_39_n_0 ;
  wire \instruction[25]_i_3_n_0 ;
  wire \instruction[25]_i_40_n_0 ;
  wire \instruction[25]_i_41_n_0 ;
  wire \instruction[25]_i_42_n_0 ;
  wire \instruction[25]_i_43_n_0 ;
  wire \instruction[25]_i_44_n_0 ;
  wire \instruction[25]_i_45_n_0 ;
  wire \instruction[25]_i_46_n_0 ;
  wire \instruction[25]_i_47_n_0 ;
  wire \instruction[25]_i_5_n_0 ;
  wire \instruction[25]_i_6_n_0 ;
  wire \instruction[25]_i_7_n_0 ;
  wire \instruction[25]_i_8_n_0 ;
  wire \instruction[25]_i_9_n_0 ;
  wire \instruction[26]_i_11_n_0 ;
  wire \instruction[26]_i_12_n_0 ;
  wire \instruction[26]_i_13_n_0 ;
  wire \instruction[26]_i_14_n_0 ;
  wire \instruction[26]_i_15_n_0 ;
  wire \instruction[26]_i_16_n_0 ;
  wire \instruction[26]_i_17_n_0 ;
  wire \instruction[26]_i_18_n_0 ;
  wire \instruction[26]_i_19_n_0 ;
  wire \instruction[26]_i_1_n_0 ;
  wire \instruction[26]_i_20_n_0 ;
  wire \instruction[26]_i_22_n_0 ;
  wire \instruction[26]_i_23_n_0 ;
  wire \instruction[26]_i_24_n_0 ;
  wire \instruction[26]_i_25_n_0 ;
  wire \instruction[26]_i_2_n_0 ;
  wire \instruction[26]_i_3_n_0 ;
  wire \instruction[26]_i_4_n_0 ;
  wire \instruction[26]_i_5_n_0 ;
  wire \instruction[26]_i_6_n_0 ;
  wire \instruction[26]_i_7_n_0 ;
  wire \instruction[26]_i_8_n_0 ;
  wire \instruction[26]_i_9_n_0 ;
  wire \instruction[27]_i_10_n_0 ;
  wire \instruction[27]_i_11_n_0 ;
  wire \instruction[27]_i_13_n_0 ;
  wire \instruction[27]_i_14_n_0 ;
  wire \instruction[27]_i_15_n_0 ;
  wire \instruction[27]_i_1_n_0 ;
  wire \instruction[27]_i_2_n_0 ;
  wire \instruction[27]_i_4_n_0 ;
  wire \instruction[27]_i_5_n_0 ;
  wire \instruction[27]_i_6_n_0 ;
  wire \instruction[27]_i_7_n_0 ;
  wire \instruction[27]_i_8_n_0 ;
  wire \instruction[27]_i_9_n_0 ;
  wire \instruction[2]_i_10_n_0 ;
  wire \instruction[2]_i_11_n_0 ;
  wire \instruction[2]_i_12_n_0 ;
  wire \instruction[2]_i_13_n_0 ;
  wire \instruction[2]_i_14_n_0 ;
  wire \instruction[2]_i_15_n_0 ;
  wire \instruction[2]_i_17_n_0 ;
  wire \instruction[2]_i_18_n_0 ;
  wire \instruction[2]_i_1_n_0 ;
  wire \instruction[2]_i_20_n_0 ;
  wire \instruction[2]_i_21_n_0 ;
  wire \instruction[2]_i_22_n_0 ;
  wire \instruction[2]_i_23_n_0 ;
  wire \instruction[2]_i_24_n_0 ;
  wire \instruction[2]_i_25_n_0 ;
  wire \instruction[2]_i_26_n_0 ;
  wire \instruction[2]_i_27_n_0 ;
  wire \instruction[2]_i_29_n_0 ;
  wire \instruction[2]_i_32_n_0 ;
  wire \instruction[2]_i_33_n_0 ;
  wire \instruction[2]_i_34_n_0 ;
  wire \instruction[2]_i_35_n_0 ;
  wire \instruction[2]_i_36_n_0 ;
  wire \instruction[2]_i_39_n_0 ;
  wire \instruction[2]_i_3_n_0 ;
  wire \instruction[2]_i_40_n_0 ;
  wire \instruction[2]_i_41_n_0 ;
  wire \instruction[2]_i_42_n_0 ;
  wire \instruction[2]_i_43_n_0 ;
  wire \instruction[2]_i_44_n_0 ;
  wire \instruction[2]_i_45_n_0 ;
  wire \instruction[2]_i_46_n_0 ;
  wire \instruction[2]_i_47_n_0 ;
  wire \instruction[2]_i_49_n_0 ;
  wire \instruction[2]_i_50_n_0 ;
  wire \instruction[2]_i_51_n_0 ;
  wire \instruction[2]_i_52_n_0 ;
  wire \instruction[2]_i_53_n_0 ;
  wire \instruction[2]_i_54_n_0 ;
  wire \instruction[2]_i_55_n_0 ;
  wire \instruction[2]_i_56_n_0 ;
  wire \instruction[2]_i_6_n_0 ;
  wire \instruction[2]_i_7_n_0 ;
  wire \instruction[2]_i_8_n_0 ;
  wire \instruction[2]_i_9_n_0 ;
  wire \instruction[3]_i_10_n_0 ;
  wire \instruction[3]_i_11_n_0 ;
  wire \instruction[3]_i_12_n_0 ;
  wire \instruction[3]_i_15_n_0 ;
  wire \instruction[3]_i_16_n_0 ;
  wire \instruction[3]_i_19_n_0 ;
  wire \instruction[3]_i_1_n_0 ;
  wire \instruction[3]_i_20_n_0 ;
  wire \instruction[3]_i_21_n_0 ;
  wire \instruction[3]_i_23_n_0 ;
  wire \instruction[3]_i_25_n_0 ;
  wire \instruction[3]_i_26_n_0 ;
  wire \instruction[3]_i_27_n_0 ;
  wire \instruction[3]_i_28_n_0 ;
  wire \instruction[3]_i_29_n_0 ;
  wire \instruction[3]_i_2_n_0 ;
  wire \instruction[3]_i_30_n_0 ;
  wire \instruction[3]_i_31_n_0 ;
  wire \instruction[3]_i_32_n_0 ;
  wire \instruction[3]_i_33_n_0 ;
  wire \instruction[3]_i_34_n_0 ;
  wire \instruction[3]_i_35_n_0 ;
  wire \instruction[3]_i_36_n_0 ;
  wire \instruction[3]_i_37_n_0 ;
  wire \instruction[3]_i_38_n_0 ;
  wire \instruction[3]_i_39_n_0 ;
  wire \instruction[3]_i_40_n_0 ;
  wire \instruction[3]_i_41_n_0 ;
  wire \instruction[3]_i_42_n_0 ;
  wire \instruction[3]_i_43_n_0 ;
  wire \instruction[3]_i_44_n_0 ;
  wire \instruction[3]_i_45_n_0 ;
  wire \instruction[3]_i_46_n_0 ;
  wire \instruction[3]_i_47_n_0 ;
  wire \instruction[3]_i_48_n_0 ;
  wire \instruction[3]_i_49_n_0 ;
  wire \instruction[3]_i_4_n_0 ;
  wire \instruction[3]_i_50_n_0 ;
  wire \instruction[3]_i_51_n_0 ;
  wire \instruction[3]_i_54_n_0 ;
  wire \instruction[3]_i_55_n_0 ;
  wire \instruction[3]_i_58_n_0 ;
  wire \instruction[3]_i_60_n_0 ;
  wire \instruction[3]_i_61_n_0 ;
  wire \instruction[3]_i_62_n_0 ;
  wire \instruction[3]_i_63_n_0 ;
  wire \instruction[3]_i_64_n_0 ;
  wire \instruction[3]_i_66_n_0 ;
  wire \instruction[3]_i_67_n_0 ;
  wire \instruction[3]_i_68_n_0 ;
  wire \instruction[3]_i_69_n_0 ;
  wire \instruction[3]_i_6_n_0 ;
  wire \instruction[3]_i_70_n_0 ;
  wire \instruction[3]_i_71_n_0 ;
  wire \instruction[3]_i_72_n_0 ;
  wire \instruction[3]_i_73_n_0 ;
  wire \instruction[3]_i_74_n_0 ;
  wire \instruction[3]_i_75_n_0 ;
  wire \instruction[3]_i_76_n_0 ;
  wire \instruction[3]_i_77_n_0 ;
  wire \instruction[3]_i_78_n_0 ;
  wire \instruction[3]_i_79_n_0 ;
  wire \instruction[3]_i_7_n_0 ;
  wire \instruction[3]_i_80_n_0 ;
  wire \instruction[3]_i_81_n_0 ;
  wire \instruction[3]_i_82_n_0 ;
  wire \instruction[3]_i_83_n_0 ;
  wire \instruction[3]_i_8_n_0 ;
  wire \instruction[3]_i_9_n_0 ;
  wire \instruction[4]_i_12_n_0 ;
  wire \instruction[4]_i_14_n_0 ;
  wire \instruction[4]_i_15_n_0 ;
  wire \instruction[4]_i_16_n_0 ;
  wire \instruction[4]_i_17_n_0 ;
  wire \instruction[4]_i_18_n_0 ;
  wire \instruction[4]_i_19_n_0 ;
  wire \instruction[4]_i_1_n_0 ;
  wire \instruction[4]_i_20_n_0 ;
  wire \instruction[4]_i_21_n_0 ;
  wire \instruction[4]_i_22_n_0 ;
  wire \instruction[4]_i_23_n_0 ;
  wire \instruction[4]_i_24_n_0 ;
  wire \instruction[4]_i_28_n_0 ;
  wire \instruction[4]_i_29_n_0 ;
  wire \instruction[4]_i_2_n_0 ;
  wire \instruction[4]_i_31_n_0 ;
  wire \instruction[4]_i_32_n_0 ;
  wire \instruction[4]_i_33_n_0 ;
  wire \instruction[4]_i_34_n_0 ;
  wire \instruction[4]_i_35_n_0 ;
  wire \instruction[4]_i_37_n_0 ;
  wire \instruction[4]_i_38_n_0 ;
  wire \instruction[4]_i_39_n_0 ;
  wire \instruction[4]_i_3_n_0 ;
  wire \instruction[4]_i_40_n_0 ;
  wire \instruction[4]_i_41_n_0 ;
  wire \instruction[4]_i_42_n_0 ;
  wire \instruction[4]_i_43_n_0 ;
  wire \instruction[4]_i_44_n_0 ;
  wire \instruction[4]_i_45_n_0 ;
  wire \instruction[4]_i_46_n_0 ;
  wire \instruction[4]_i_47_n_0 ;
  wire \instruction[4]_i_48_n_0 ;
  wire \instruction[4]_i_50_n_0 ;
  wire \instruction[4]_i_51_n_0 ;
  wire \instruction[4]_i_5_n_0 ;
  wire \instruction[4]_i_7_n_0 ;
  wire \instruction[4]_i_8_n_0 ;
  wire \instruction[4]_i_9_n_0 ;
  wire \instruction[5]_i_10_n_0 ;
  wire \instruction[5]_i_11_n_0 ;
  wire \instruction[5]_i_12_n_0 ;
  wire \instruction[5]_i_13_n_0 ;
  wire \instruction[5]_i_14_n_0 ;
  wire \instruction[5]_i_17_n_0 ;
  wire \instruction[5]_i_1_n_0 ;
  wire \instruction[5]_i_20_n_0 ;
  wire \instruction[5]_i_21_n_0 ;
  wire \instruction[5]_i_22_n_0 ;
  wire \instruction[5]_i_24_n_0 ;
  wire \instruction[5]_i_25_n_0 ;
  wire \instruction[5]_i_26_n_0 ;
  wire \instruction[5]_i_27_n_0 ;
  wire \instruction[5]_i_28_n_0 ;
  wire \instruction[5]_i_29_n_0 ;
  wire \instruction[5]_i_2_n_0 ;
  wire \instruction[5]_i_30_n_0 ;
  wire \instruction[5]_i_31_n_0 ;
  wire \instruction[5]_i_32_n_0 ;
  wire \instruction[5]_i_33_n_0 ;
  wire \instruction[5]_i_34_n_0 ;
  wire \instruction[5]_i_37_n_0 ;
  wire \instruction[5]_i_39_n_0 ;
  wire \instruction[5]_i_3_n_0 ;
  wire \instruction[5]_i_42_n_0 ;
  wire \instruction[5]_i_43_n_0 ;
  wire \instruction[5]_i_44_n_0 ;
  wire \instruction[5]_i_45_n_0 ;
  wire \instruction[5]_i_46_n_0 ;
  wire \instruction[5]_i_47_n_0 ;
  wire \instruction[5]_i_48_n_0 ;
  wire \instruction[5]_i_49_n_0 ;
  wire \instruction[5]_i_6_n_0 ;
  wire \instruction[5]_i_7_n_0 ;
  wire \instruction[5]_i_8_n_0 ;
  wire \instruction[5]_i_9_n_0 ;
  wire \instruction[6]_i_10_n_0 ;
  wire \instruction[6]_i_12_n_0 ;
  wire \instruction[6]_i_13_n_0 ;
  wire \instruction[6]_i_14_n_0 ;
  wire \instruction[6]_i_15_n_0 ;
  wire \instruction[6]_i_16_n_0 ;
  wire \instruction[6]_i_17_n_0 ;
  wire \instruction[6]_i_18_n_0 ;
  wire \instruction[6]_i_19_n_0 ;
  wire \instruction[6]_i_1_n_0 ;
  wire \instruction[6]_i_20_n_0 ;
  wire \instruction[6]_i_23_n_0 ;
  wire \instruction[6]_i_24_n_0 ;
  wire \instruction[6]_i_25_n_0 ;
  wire \instruction[6]_i_26_n_0 ;
  wire \instruction[6]_i_28_n_0 ;
  wire \instruction[6]_i_31_n_0 ;
  wire \instruction[6]_i_33_n_0 ;
  wire \instruction[6]_i_34_n_0 ;
  wire \instruction[6]_i_35_n_0 ;
  wire \instruction[6]_i_36_n_0 ;
  wire \instruction[6]_i_38_n_0 ;
  wire \instruction[6]_i_39_n_0 ;
  wire \instruction[6]_i_3_n_0 ;
  wire \instruction[6]_i_40_n_0 ;
  wire \instruction[6]_i_41_n_0 ;
  wire \instruction[6]_i_42_n_0 ;
  wire \instruction[6]_i_43_n_0 ;
  wire \instruction[6]_i_44_n_0 ;
  wire \instruction[6]_i_45_n_0 ;
  wire \instruction[6]_i_46_n_0 ;
  wire \instruction[6]_i_47_n_0 ;
  wire \instruction[6]_i_48_n_0 ;
  wire \instruction[6]_i_49_n_0 ;
  wire \instruction[6]_i_4_n_0 ;
  wire \instruction[6]_i_50_n_0 ;
  wire \instruction[6]_i_51_n_0 ;
  wire \instruction[6]_i_5_n_0 ;
  wire \instruction[6]_i_9_n_0 ;
  wire \instruction[7]_i_10_n_0 ;
  wire \instruction[7]_i_11_n_0 ;
  wire \instruction[7]_i_12_n_0 ;
  wire \instruction[7]_i_13_n_0 ;
  wire \instruction[7]_i_14_n_0 ;
  wire \instruction[7]_i_16_n_0 ;
  wire \instruction[7]_i_17_n_0 ;
  wire \instruction[7]_i_18_n_0 ;
  wire \instruction[7]_i_19_n_0 ;
  wire \instruction[7]_i_1_n_0 ;
  wire \instruction[7]_i_20_n_0 ;
  wire \instruction[7]_i_21_n_0 ;
  wire \instruction[7]_i_22_n_0 ;
  wire \instruction[7]_i_23_n_0 ;
  wire \instruction[7]_i_24_n_0 ;
  wire \instruction[7]_i_25_n_0 ;
  wire \instruction[7]_i_26_n_0 ;
  wire \instruction[7]_i_27_n_0 ;
  wire \instruction[7]_i_28_n_0 ;
  wire \instruction[7]_i_29_n_0 ;
  wire \instruction[7]_i_2_n_0 ;
  wire \instruction[7]_i_30_n_0 ;
  wire \instruction[7]_i_3_n_0 ;
  wire \instruction[7]_i_4_n_0 ;
  wire \instruction[7]_i_5_n_0 ;
  wire \instruction[7]_i_6_n_0 ;
  wire \instruction[7]_i_7_n_0 ;
  wire \instruction[7]_i_8_n_0 ;
  wire \instruction[8]_i_10_n_0 ;
  wire \instruction[8]_i_11_n_0 ;
  wire \instruction[8]_i_12_n_0 ;
  wire \instruction[8]_i_13_n_0 ;
  wire \instruction[8]_i_1_n_0 ;
  wire \instruction[8]_i_3_n_0 ;
  wire \instruction[8]_i_4_n_0 ;
  wire \instruction[8]_i_5_n_0 ;
  wire \instruction[8]_i_6_n_0 ;
  wire \instruction[8]_i_7_n_0 ;
  wire \instruction[8]_i_8_n_0 ;
  wire \instruction[9]_i_10_n_0 ;
  wire \instruction[9]_i_11_n_0 ;
  wire \instruction[9]_i_12_n_0 ;
  wire \instruction[9]_i_13_n_0 ;
  wire \instruction[9]_i_14_n_0 ;
  wire \instruction[9]_i_1_n_0 ;
  wire \instruction[9]_i_2_n_0 ;
  wire \instruction[9]_i_3_n_0 ;
  wire \instruction[9]_i_4_n_0 ;
  wire \instruction[9]_i_6_n_0 ;
  wire \instruction[9]_i_7_n_0 ;
  wire \instruction[9]_i_8_n_0 ;
  wire \instruction[9]_i_9_n_0 ;
  wire \instruction_reg[0]_i_10_n_0 ;
  wire \instruction_reg[0]_i_20_n_0 ;
  wire \instruction_reg[0]_i_24_n_0 ;
  wire \instruction_reg[0]_i_27_n_0 ;
  wire \instruction_reg[0]_i_2_n_0 ;
  wire \instruction_reg[0]_i_33_n_0 ;
  wire \instruction_reg[0]_i_36_n_0 ;
  wire \instruction_reg[0]_i_37_n_0 ;
  wire \instruction_reg[0]_i_39_n_0 ;
  wire \instruction_reg[0]_i_47_n_0 ;
  wire \instruction_reg[0]_i_4_n_0 ;
  wire \instruction_reg[0]_i_50_n_0 ;
  wire \instruction_reg[0]_i_5_n_0 ;
  wire \instruction_reg[16]_i_17_n_0 ;
  wire \instruction_reg[16]_i_18_n_0 ;
  wire \instruction_reg[16]_i_22_n_0 ;
  wire \instruction_reg[16]_i_3_n_0 ;
  wire \instruction_reg[16]_i_5_n_0 ;
  wire \instruction_reg[17]_i_12_n_0 ;
  wire \instruction_reg[17]_i_14_n_0 ;
  wire \instruction_reg[17]_i_26_n_0 ;
  wire \instruction_reg[17]_i_30_n_0 ;
  wire \instruction_reg[17]_i_3_n_0 ;
  wire \instruction_reg[17]_i_46_n_0 ;
  wire \instruction_reg[17]_i_4_n_0 ;
  wire \instruction_reg[18]_i_10_n_0 ;
  wire \instruction_reg[18]_i_12_n_0 ;
  wire \instruction_reg[18]_i_13_n_0 ;
  wire \instruction_reg[18]_i_21_n_0 ;
  wire \instruction_reg[18]_i_22_n_0 ;
  wire \instruction_reg[18]_i_23_n_0 ;
  wire \instruction_reg[18]_i_4_n_0 ;
  wire \instruction_reg[18]_i_5_n_0 ;
  wire \instruction_reg[18]_i_8_n_0 ;
  wire \instruction_reg[19]_i_10_n_0 ;
  wire \instruction_reg[19]_i_12_n_0 ;
  wire \instruction_reg[1]_i_17_n_0 ;
  wire \instruction_reg[1]_i_18_n_0 ;
  wire \instruction_reg[1]_i_23_n_0 ;
  wire \instruction_reg[1]_i_24_n_0 ;
  wire \instruction_reg[1]_i_2_n_0 ;
  wire \instruction_reg[1]_i_48_n_0 ;
  wire \instruction_reg[1]_i_4_n_0 ;
  wire \instruction_reg[1]_i_50_n_0 ;
  wire \instruction_reg[1]_i_52_n_0 ;
  wire \instruction_reg[1]_i_53_n_0 ;
  wire \instruction_reg[1]_i_5_n_0 ;
  wire \instruction_reg[1]_i_6_n_0 ;
  wire \instruction_reg[1]_i_7_n_0 ;
  wire \instruction_reg[20]_i_12_n_0 ;
  wire \instruction_reg[20]_i_23_n_0 ;
  wire \instruction_reg[20]_i_25_n_0 ;
  wire \instruction_reg[20]_i_8_n_0 ;
  wire \instruction_reg[21]_i_10_n_0 ;
  wire \instruction_reg[21]_i_11_n_0 ;
  wire \instruction_reg[21]_i_13_n_0 ;
  wire \instruction_reg[21]_i_33_n_0 ;
  wire \instruction_reg[21]_i_34_n_0 ;
  wire \instruction_reg[21]_i_35_n_0 ;
  wire \instruction_reg[21]_i_36_n_0 ;
  wire \instruction_reg[21]_i_39_n_0 ;
  wire \instruction_reg[21]_i_40_n_0 ;
  wire \instruction_reg[21]_i_44_n_0 ;
  wire \instruction_reg[21]_i_4_n_0 ;
  wire \instruction_reg[21]_i_5_n_0 ;
  wire \instruction_reg[22]_i_5_n_0 ;
  wire \instruction_reg[23]_i_10_n_0 ;
  wire \instruction_reg[23]_i_27_n_0 ;
  wire \instruction_reg[23]_i_2_n_0 ;
  wire \instruction_reg[23]_i_33_n_0 ;
  wire \instruction_reg[23]_i_40_n_0 ;
  wire \instruction_reg[23]_i_43_n_0 ;
  wire \instruction_reg[23]_i_44_n_0 ;
  wire \instruction_reg[23]_i_45_n_0 ;
  wire \instruction_reg[23]_i_4_n_0 ;
  wire \instruction_reg[23]_i_5_n_0 ;
  wire \instruction_reg[23]_i_6_n_0 ;
  wire \instruction_reg[24]_i_19_n_0 ;
  wire \instruction_reg[24]_i_20_n_0 ;
  wire \instruction_reg[24]_i_25_n_0 ;
  wire \instruction_reg[24]_i_3_n_0 ;
  wire \instruction_reg[24]_i_41_n_0 ;
  wire \instruction_reg[24]_i_45_n_0 ;
  wire \instruction_reg[24]_i_4_n_0 ;
  wire \instruction_reg[24]_i_5_n_0 ;
  wire \instruction_reg[25]_i_19_n_0 ;
  wire \instruction_reg[25]_i_20_n_0 ;
  wire \instruction_reg[25]_i_26_n_0 ;
  wire \instruction_reg[25]_i_31_n_0 ;
  wire \instruction_reg[25]_i_32_n_0 ;
  wire \instruction_reg[25]_i_33_n_0 ;
  wire \instruction_reg[25]_i_34_n_0 ;
  wire \instruction_reg[25]_i_4_n_0 ;
  wire \instruction_reg[26]_i_10_n_0 ;
  wire \instruction_reg[26]_i_21_n_0 ;
  wire \instruction_reg[27]_i_12_n_0 ;
  wire \instruction_reg[27]_i_3_n_0 ;
  wire \instruction_reg[2]_i_16_n_0 ;
  wire \instruction_reg[2]_i_19_n_0 ;
  wire \instruction_reg[2]_i_28_n_0 ;
  wire \instruction_reg[2]_i_2_n_0 ;
  wire \instruction_reg[2]_i_30_n_0 ;
  wire \instruction_reg[2]_i_31_n_0 ;
  wire \instruction_reg[2]_i_37_n_0 ;
  wire \instruction_reg[2]_i_38_n_0 ;
  wire \instruction_reg[2]_i_48_n_0 ;
  wire \instruction_reg[2]_i_4_n_0 ;
  wire \instruction_reg[2]_i_5_n_0 ;
  wire \instruction_reg[3]_i_13_n_0 ;
  wire \instruction_reg[3]_i_14_n_0 ;
  wire \instruction_reg[3]_i_17_n_0 ;
  wire \instruction_reg[3]_i_18_n_0 ;
  wire \instruction_reg[3]_i_22_n_0 ;
  wire \instruction_reg[3]_i_24_n_0 ;
  wire \instruction_reg[3]_i_3_n_0 ;
  wire \instruction_reg[3]_i_52_n_0 ;
  wire \instruction_reg[3]_i_53_n_0 ;
  wire \instruction_reg[3]_i_56_n_0 ;
  wire \instruction_reg[3]_i_57_n_0 ;
  wire \instruction_reg[3]_i_59_n_0 ;
  wire \instruction_reg[3]_i_5_n_0 ;
  wire \instruction_reg[3]_i_65_n_0 ;
  wire \instruction_reg[4]_i_10_n_0 ;
  wire \instruction_reg[4]_i_11_n_0 ;
  wire \instruction_reg[4]_i_13_n_0 ;
  wire \instruction_reg[4]_i_25_n_0 ;
  wire \instruction_reg[4]_i_26_n_0 ;
  wire \instruction_reg[4]_i_27_n_0 ;
  wire \instruction_reg[4]_i_30_n_0 ;
  wire \instruction_reg[4]_i_36_n_0 ;
  wire \instruction_reg[4]_i_49_n_0 ;
  wire \instruction_reg[4]_i_4_n_0 ;
  wire \instruction_reg[4]_i_6_n_0 ;
  wire \instruction_reg[5]_i_15_n_0 ;
  wire \instruction_reg[5]_i_16_n_0 ;
  wire \instruction_reg[5]_i_18_n_0 ;
  wire \instruction_reg[5]_i_19_n_0 ;
  wire \instruction_reg[5]_i_23_n_0 ;
  wire \instruction_reg[5]_i_35_n_0 ;
  wire \instruction_reg[5]_i_36_n_0 ;
  wire \instruction_reg[5]_i_38_n_0 ;
  wire \instruction_reg[5]_i_40_n_0 ;
  wire \instruction_reg[5]_i_41_n_0 ;
  wire \instruction_reg[5]_i_4_n_0 ;
  wire \instruction_reg[5]_i_5_n_0 ;
  wire \instruction_reg[6]_i_11_n_0 ;
  wire \instruction_reg[6]_i_21_n_0 ;
  wire \instruction_reg[6]_i_22_n_0 ;
  wire \instruction_reg[6]_i_27_n_0 ;
  wire \instruction_reg[6]_i_29_n_0 ;
  wire \instruction_reg[6]_i_2_n_0 ;
  wire \instruction_reg[6]_i_30_n_0 ;
  wire \instruction_reg[6]_i_32_n_0 ;
  wire \instruction_reg[6]_i_37_n_0 ;
  wire \instruction_reg[6]_i_6_n_0 ;
  wire \instruction_reg[6]_i_7_n_0 ;
  wire \instruction_reg[6]_i_8_n_0 ;
  wire \instruction_reg[7]_i_15_n_0 ;
  wire \instruction_reg[7]_i_9_n_0 ;
  wire \instruction_reg[8]_i_2_n_0 ;
  wire \instruction_reg[8]_i_9_n_0 ;
  wire \instruction_reg[9]_i_5_n_0 ;
  wire \instruction_reg_n_0_[0] ;
  wire \instruction_reg_n_0_[15] ;
  wire \instruction_reg_n_0_[1] ;
  wire \instruction_reg_n_0_[2] ;
  wire \instruction_reg_n_0_[3] ;
  wire \instruction_reg_n_0_[4] ;
  wire \instruction_reg_n_0_[5] ;
  wire \instruction_reg_n_0_[6] ;
  wire \instruction_reg_n_0_[7] ;
  wire \instruction_reg_n_0_[8] ;
  wire \instruction_reg_n_0_[9] ;
  wire [15:4]literal_2;
  wire [31:0]load_data;
  wire memory_reg_0_i_2_n_0;
  wire memory_reg_1_ENARDEN_cooolgate_en_sig_1;
  wire memory_reg_2_ENARDEN_cooolgate_en_sig_2;
  wire memory_reg_3_ENARDEN_cooolgate_en_sig_3;
  wire memory_reg_4_ENARDEN_cooolgate_en_sig_4;
  wire memory_reg_5_ENARDEN_cooolgate_en_sig_5;
  wire memory_reg_6_ENARDEN_cooolgate_en_sig_6;
  wire memory_reg_7_ENARDEN_cooolgate_en_sig_7;
  wire [3:0]opcode;
  wire [3:0]opcode_2;
  wire opcode_20;
  wire operand_a1;
  wire operand_b1;
  wire p_0_in;
  wire \program_counter[10]_i_1_n_0 ;
  wire \program_counter[11]_i_1_n_0 ;
  wire \program_counter[12]_i_1_n_0 ;
  wire \program_counter[13]_i_1_n_0 ;
  wire \program_counter[14]_i_1_n_0 ;
  wire \program_counter[15]_i_11_n_0 ;
  wire \program_counter[15]_i_12_n_0 ;
  wire \program_counter[15]_i_13_n_0 ;
  wire \program_counter[15]_i_14_n_0 ;
  wire \program_counter[15]_i_15_n_0 ;
  wire \program_counter[15]_i_16_n_0 ;
  wire \program_counter[15]_i_17_n_0 ;
  wire \program_counter[15]_i_18_n_0 ;
  wire \program_counter[15]_i_1_n_0 ;
  wire \program_counter[15]_i_2_n_0 ;
  wire \program_counter[15]_i_4_n_0 ;
  wire \program_counter[15]_i_5_n_0 ;
  wire \program_counter[15]_i_6_n_0 ;
  wire \program_counter[15]_i_7_n_0 ;
  wire [15:0]program_counter_1;
  wire [15:0]program_counter_2;
  wire \program_counter_reg_n_0_[0] ;
  wire \program_counter_reg_n_0_[10] ;
  wire \program_counter_reg_n_0_[11] ;
  wire \program_counter_reg_n_0_[12] ;
  wire \program_counter_reg_n_0_[13] ;
  wire \program_counter_reg_n_0_[14] ;
  wire \program_counter_reg_n_0_[15] ;
  wire \program_counter_reg_n_0_[1] ;
  wire \program_counter_reg_n_0_[2] ;
  wire \program_counter_reg_n_0_[3] ;
  wire \program_counter_reg_n_0_[4] ;
  wire \program_counter_reg_n_0_[5] ;
  wire \program_counter_reg_n_0_[6] ;
  wire \program_counter_reg_n_0_[7] ;
  wire \program_counter_reg_n_0_[8] ;
  wire \program_counter_reg_n_0_[9] ;
  wire \program_counter_reg_rep[2]_rep__0_n_0 ;
  wire \program_counter_reg_rep[2]_rep_n_0 ;
  wire \program_counter_reg_rep[3]_rep__0_n_0 ;
  wire \program_counter_reg_rep[3]_rep__1_n_0 ;
  wire \program_counter_reg_rep[3]_rep_n_0 ;
  wire \program_counter_reg_rep[4]_i_2_n_0 ;
  wire \program_counter_reg_rep[4]_rep__0_n_0 ;
  wire \program_counter_reg_rep[4]_rep__1_n_0 ;
  wire \program_counter_reg_rep[4]_rep__2_n_0 ;
  wire \program_counter_reg_rep[4]_rep_n_0 ;
  wire \program_counter_reg_rep[5]_rep__0_n_0 ;
  wire \program_counter_reg_rep[5]_rep__1_n_0 ;
  wire \program_counter_reg_rep[5]_rep__2_n_0 ;
  wire \program_counter_reg_rep[5]_rep_n_0 ;
  wire \program_counter_reg_rep[6]_rep__0_n_0 ;
  wire \program_counter_reg_rep[6]_rep__1_n_0 ;
  wire \program_counter_reg_rep[6]_rep__2_n_0 ;
  wire \program_counter_reg_rep[6]_rep_n_0 ;
  wire \program_counter_reg_rep[7]_rep__0_n_0 ;
  wire \program_counter_reg_rep[7]_rep__1_n_0 ;
  wire \program_counter_reg_rep[7]_rep_n_0 ;
  wire \program_counter_reg_rep[8]_i_2_n_0 ;
  wire \program_counter_reg_rep[8]_rep__0_n_0 ;
  wire \program_counter_reg_rep[8]_rep__1_n_0 ;
  wire \program_counter_reg_rep[8]_rep__2_n_0 ;
  wire \program_counter_reg_rep[8]_rep_n_0 ;
  wire \program_counter_reg_rep[9]_i_5_n_0 ;
  wire \program_counter_reg_rep[9]_rep__0_n_0 ;
  wire \program_counter_reg_rep[9]_rep__1_n_0 ;
  wire \program_counter_reg_rep[9]_rep__2_n_0 ;
  wire \program_counter_reg_rep[9]_rep_n_0 ;
  wire \program_counter_reg_rep_n_0_[0] ;
  wire \program_counter_reg_rep_n_0_[1] ;
  wire \program_counter_reg_rep_n_0_[2] ;
  wire \program_counter_reg_rep_n_0_[3] ;
  wire \program_counter_reg_rep_n_0_[4] ;
  wire \program_counter_reg_rep_n_0_[5] ;
  wire \program_counter_reg_rep_n_0_[6] ;
  wire \program_counter_reg_rep_n_0_[7] ;
  wire \program_counter_reg_rep_n_0_[8] ;
  wire \program_counter_reg_rep_n_0_[9] ;
  wire \program_counter_rep[0]_i_1_n_0 ;
  wire \program_counter_rep[1]_i_1_n_0 ;
  wire \program_counter_rep[2]_i_1_n_0 ;
  wire \program_counter_rep[3]_i_1_n_0 ;
  wire \program_counter_rep[4]_i_1_n_0 ;
  wire \program_counter_rep[5]_i_1_n_0 ;
  wire \program_counter_rep[6]_i_1_n_0 ;
  wire \program_counter_rep[7]_i_1_n_0 ;
  wire \program_counter_rep[8]_i_1_n_0 ;
  wire \program_counter_rep[9]_i_14_n_0 ;
  wire \program_counter_rep[9]_i_15_n_0 ;
  wire \program_counter_rep[9]_i_16_n_0 ;
  wire \program_counter_rep[9]_i_17_n_0 ;
  wire \program_counter_rep[9]_i_18_n_0 ;
  wire \program_counter_rep[9]_i_19_n_0 ;
  wire \program_counter_rep[9]_i_20_n_0 ;
  wire \program_counter_rep[9]_i_21_n_0 ;
  wire \program_counter_rep[9]_i_22_n_0 ;
  wire \program_counter_rep[9]_i_2_n_0 ;
  wire \program_counter_rep[9]_i_3_n_0 ;
  wire \program_counter_rep[9]_i_4_n_0 ;
  wire \program_counter_rep[9]_i_6_n_0 ;
  wire \program_counter_rep[9]_i_7_n_0 ;
  wire \program_counter_rep[9]_i_8_n_0 ;
  wire \program_counter_rep[9]_i_9_n_0 ;
  wire [31:0]read_input;
  wire \read_input[31]_i_1_n_0 ;
  wire \read_input[31]_i_2_n_0 ;
  wire [31:0]register_a;
  wire [31:0]register_b;
  wire [31:0]result;
  wire \result[0]_i_10_n_0 ;
  wire \result[0]_i_12_n_0 ;
  wire \result[0]_i_13_n_0 ;
  wire \result[0]_i_14_n_0 ;
  wire \result[0]_i_15_n_0 ;
  wire \result[0]_i_16_n_0 ;
  wire \result[0]_i_17_n_0 ;
  wire \result[0]_i_18_n_0 ;
  wire \result[0]_i_19_n_0 ;
  wire \result[0]_i_1_n_0 ;
  wire \result[0]_i_2_n_0 ;
  wire \result[0]_i_3_n_0 ;
  wire \result[0]_i_5_n_0 ;
  wire \result[0]_i_6_n_0 ;
  wire \result[0]_i_8_n_0 ;
  wire \result[0]_i_9_n_0 ;
  wire \result[10]_i_1_n_0 ;
  wire \result[10]_i_2_n_0 ;
  wire \result[11]_i_10_n_0 ;
  wire \result[11]_i_11_n_0 ;
  wire \result[11]_i_12_n_0 ;
  wire \result[11]_i_13_n_0 ;
  wire \result[11]_i_14_n_0 ;
  wire \result[11]_i_15_n_0 ;
  wire \result[11]_i_16_n_0 ;
  wire \result[11]_i_17_n_0 ;
  wire \result[11]_i_18_n_0 ;
  wire \result[11]_i_1_n_0 ;
  wire \result[11]_i_2_n_0 ;
  wire \result[11]_i_3_n_0 ;
  wire \result[11]_i_7_n_0 ;
  wire \result[11]_i_8_n_0 ;
  wire \result[11]_i_9_n_0 ;
  wire \result[12]_i_1_n_0 ;
  wire \result[12]_i_2_n_0 ;
  wire \result[12]_i_4_n_0 ;
  wire \result[13]_i_1_n_0 ;
  wire \result[13]_i_2_n_0 ;
  wire \result[13]_i_3_n_0 ;
  wire \result[14]_i_1_n_0 ;
  wire \result[14]_i_2_n_0 ;
  wire \result[14]_i_3_n_0 ;
  wire \result[15]_i_1_n_0 ;
  wire \result[15]_i_3_n_0 ;
  wire \result[15]_i_4_n_0 ;
  wire \result[15]_i_5_n_0 ;
  wire \result[15]_i_6_n_0 ;
  wire \result[15]_i_7_n_0 ;
  wire \result[15]_i_8_n_0 ;
  wire \result[16]_i_10_n_0 ;
  wire \result[16]_i_11_n_0 ;
  wire \result[16]_i_12_n_0 ;
  wire \result[16]_i_13_n_0 ;
  wire \result[16]_i_14_n_0 ;
  wire \result[16]_i_15_n_0 ;
  wire \result[16]_i_16_n_0 ;
  wire \result[16]_i_17_n_0 ;
  wire \result[16]_i_1_n_0 ;
  wire \result[16]_i_21_n_0 ;
  wire \result[16]_i_22_n_0 ;
  wire \result[16]_i_23_n_0 ;
  wire \result[16]_i_24_n_0 ;
  wire \result[16]_i_2_n_0 ;
  wire \result[16]_i_3_n_0 ;
  wire \result[16]_i_5_n_0 ;
  wire \result[16]_i_7_n_0 ;
  wire \result[17]_i_1_n_0 ;
  wire \result[17]_i_2_n_0 ;
  wire \result[18]_i_1_n_0 ;
  wire \result[18]_i_2_n_0 ;
  wire \result[19]_i_10_n_0 ;
  wire \result[19]_i_11_n_0 ;
  wire \result[19]_i_12_n_0 ;
  wire \result[19]_i_1_n_0 ;
  wire \result[19]_i_3_n_0 ;
  wire \result[19]_i_5_n_0 ;
  wire \result[19]_i_6_n_0 ;
  wire \result[19]_i_7_n_0 ;
  wire \result[19]_i_8_n_0 ;
  wire \result[19]_i_9_n_0 ;
  wire \result[1]_i_1_n_0 ;
  wire \result[1]_i_2_n_0 ;
  wire \result[1]_i_3_n_0 ;
  wire \result[1]_i_4_n_0 ;
  wire \result[20]_i_1_n_0 ;
  wire \result[20]_i_2_n_0 ;
  wire \result[21]_i_1_n_0 ;
  wire \result[21]_i_2_n_0 ;
  wire \result[22]_i_1_n_0 ;
  wire \result[22]_i_2_n_0 ;
  wire \result[23]_i_10_n_0 ;
  wire \result[23]_i_11_n_0 ;
  wire \result[23]_i_12_n_0 ;
  wire \result[23]_i_13_n_0 ;
  wire \result[23]_i_14_n_0 ;
  wire \result[23]_i_15_n_0 ;
  wire \result[23]_i_16_n_0 ;
  wire \result[23]_i_17_n_0 ;
  wire \result[23]_i_1_n_0 ;
  wire \result[23]_i_3_n_0 ;
  wire \result[23]_i_4_n_0 ;
  wire \result[23]_i_5_n_0 ;
  wire \result[23]_i_6_n_0 ;
  wire \result[23]_i_7_n_0 ;
  wire \result[24]_i_1_n_0 ;
  wire \result[24]_i_2_n_0 ;
  wire \result[25]_i_1_n_0 ;
  wire \result[25]_i_2_n_0 ;
  wire \result[26]_i_1_n_0 ;
  wire \result[26]_i_2_n_0 ;
  wire \result[27]_i_10_n_0 ;
  wire \result[27]_i_11_n_0 ;
  wire \result[27]_i_12_n_0 ;
  wire \result[27]_i_13_n_0 ;
  wire \result[27]_i_14_n_0 ;
  wire \result[27]_i_15_n_0 ;
  wire \result[27]_i_16_n_0 ;
  wire \result[27]_i_17_n_0 ;
  wire \result[27]_i_1_n_0 ;
  wire \result[27]_i_3_n_0 ;
  wire \result[27]_i_4_n_0 ;
  wire \result[27]_i_5_n_0 ;
  wire \result[27]_i_6_n_0 ;
  wire \result[27]_i_7_n_0 ;
  wire \result[28]_i_1_n_0 ;
  wire \result[28]_i_2_n_0 ;
  wire \result[29]_i_1_n_0 ;
  wire \result[29]_i_2_n_0 ;
  wire \result[2]_i_1_n_0 ;
  wire \result[2]_i_2_n_0 ;
  wire \result[2]_i_3_n_0 ;
  wire \result[2]_i_4_n_0 ;
  wire \result[30]_i_1_n_0 ;
  wire \result[30]_i_2_n_0 ;
  wire \result[31]_i_10_n_0 ;
  wire \result[31]_i_11_n_0 ;
  wire \result[31]_i_12_n_0 ;
  wire \result[31]_i_13_n_0 ;
  wire \result[31]_i_14_n_0 ;
  wire \result[31]_i_15_n_0 ;
  wire \result[31]_i_18_n_0 ;
  wire \result[31]_i_19_n_0 ;
  wire \result[31]_i_1_n_0 ;
  wire \result[31]_i_20_n_0 ;
  wire \result[31]_i_21_n_0 ;
  wire \result[31]_i_22_n_0 ;
  wire \result[31]_i_24_n_0 ;
  wire \result[31]_i_25_n_0 ;
  wire \result[31]_i_26_n_0 ;
  wire \result[31]_i_27_n_0 ;
  wire \result[31]_i_28_n_0 ;
  wire \result[31]_i_29_n_0 ;
  wire \result[31]_i_2_n_0 ;
  wire \result[31]_i_30_n_0 ;
  wire \result[31]_i_31_n_0 ;
  wire \result[31]_i_3_n_0 ;
  wire \result[31]_i_6_n_0 ;
  wire \result[31]_i_7_n_0 ;
  wire \result[31]_i_9_n_0 ;
  wire \result[3]_i_10_n_0 ;
  wire \result[3]_i_11_n_0 ;
  wire \result[3]_i_12_n_0 ;
  wire \result[3]_i_13_n_0 ;
  wire \result[3]_i_14_n_0 ;
  wire \result[3]_i_15_n_0 ;
  wire \result[3]_i_16_n_0 ;
  wire \result[3]_i_17_n_0 ;
  wire \result[3]_i_18_n_0 ;
  wire \result[3]_i_19_n_0 ;
  wire \result[3]_i_1_n_0 ;
  wire \result[3]_i_2_n_0 ;
  wire \result[3]_i_4_n_0 ;
  wire \result[3]_i_7_n_0 ;
  wire \result[3]_i_8_n_0 ;
  wire \result[3]_i_9_n_0 ;
  wire \result[4]_i_1_n_0 ;
  wire \result[4]_i_2_n_0 ;
  wire \result[4]_i_3_n_0 ;
  wire \result[4]_i_5_n_0 ;
  wire \result[5]_i_1_n_0 ;
  wire \result[5]_i_2_n_0 ;
  wire \result[5]_i_3_n_0 ;
  wire \result[5]_i_4_n_0 ;
  wire \result[6]_i_1_n_0 ;
  wire \result[6]_i_2_n_0 ;
  wire \result[6]_i_3_n_0 ;
  wire \result[6]_i_4_n_0 ;
  wire \result[7]_i_10_n_0 ;
  wire \result[7]_i_11_n_0 ;
  wire \result[7]_i_12_n_0 ;
  wire \result[7]_i_13_n_0 ;
  wire \result[7]_i_14_n_0 ;
  wire \result[7]_i_15_n_0 ;
  wire \result[7]_i_1_n_0 ;
  wire \result[7]_i_2_n_0 ;
  wire \result[7]_i_4_n_0 ;
  wire \result[7]_i_5_n_0 ;
  wire \result[7]_i_7_n_0 ;
  wire \result[7]_i_8_n_0 ;
  wire \result[7]_i_9_n_0 ;
  wire \result[8]_i_1_n_0 ;
  wire \result[8]_i_2_n_0 ;
  wire \result[8]_i_3_n_0 ;
  wire \result[9]_i_1_n_0 ;
  wire \result[9]_i_3_n_0 ;
  wire \result[9]_i_4_n_0 ;
  wire \result[9]_i_5_n_0 ;
  wire \result[9]_i_6_n_0 ;
  wire \result[9]_i_7_n_0 ;
  wire \result[9]_i_8_n_0 ;
  wire \result[9]_i_9_n_0 ;
  wire \result_reg[0]_i_11_n_0 ;
  wire \result_reg[0]_i_4_n_1 ;
  wire \result_reg[0]_i_7_n_0 ;
  wire \result_reg[11]_i_4_n_0 ;
  wire \result_reg[11]_i_5_n_0 ;
  wire \result_reg[11]_i_5_n_4 ;
  wire \result_reg[11]_i_5_n_5 ;
  wire \result_reg[11]_i_5_n_6 ;
  wire \result_reg[11]_i_5_n_7 ;
  wire \result_reg[11]_i_6_n_0 ;
  wire \result_reg[12]_i_3_n_0 ;
  wire \result_reg[15]_i_2_n_0 ;
  wire \result_reg[16]_i_4_n_0 ;
  wire \result_reg[16]_i_4_n_4 ;
  wire \result_reg[16]_i_4_n_5 ;
  wire \result_reg[16]_i_4_n_6 ;
  wire \result_reg[16]_i_4_n_7 ;
  wire \result_reg[16]_i_6_n_0 ;
  wire \result_reg[16]_i_9_n_0 ;
  wire \result_reg[16]_i_9_n_4 ;
  wire \result_reg[16]_i_9_n_5 ;
  wire \result_reg[16]_i_9_n_6 ;
  wire \result_reg[16]_i_9_n_7 ;
  wire \result_reg[19]_i_2_n_0 ;
  wire \result_reg[19]_i_4_n_0 ;
  wire \result_reg[23]_i_2_n_0 ;
  wire \result_reg[23]_i_8_n_0 ;
  wire \result_reg[23]_i_9_n_0 ;
  wire \result_reg[23]_i_9_n_4 ;
  wire \result_reg[23]_i_9_n_5 ;
  wire \result_reg[23]_i_9_n_6 ;
  wire \result_reg[23]_i_9_n_7 ;
  wire \result_reg[27]_i_2_n_0 ;
  wire \result_reg[27]_i_8_n_0 ;
  wire \result_reg[27]_i_9_n_0 ;
  wire \result_reg[27]_i_9_n_4 ;
  wire \result_reg[27]_i_9_n_5 ;
  wire \result_reg[27]_i_9_n_6 ;
  wire \result_reg[27]_i_9_n_7 ;
  wire \result_reg[31]_i_17_n_4 ;
  wire \result_reg[31]_i_17_n_5 ;
  wire \result_reg[31]_i_17_n_6 ;
  wire \result_reg[31]_i_17_n_7 ;
  wire \result_reg[3]_i_3_n_0 ;
  wire \result_reg[3]_i_3_n_4 ;
  wire \result_reg[3]_i_3_n_5 ;
  wire \result_reg[3]_i_3_n_6 ;
  wire \result_reg[3]_i_3_n_7 ;
  wire \result_reg[3]_i_5_n_0 ;
  wire \result_reg[3]_i_6_n_0 ;
  wire \result_reg[4]_i_4_n_0 ;
  wire \result_reg[7]_i_3_n_0 ;
  wire \result_reg[7]_i_3_n_4 ;
  wire \result_reg[7]_i_3_n_5 ;
  wire \result_reg[7]_i_3_n_6 ;
  wire \result_reg[7]_i_3_n_7 ;
  wire \result_reg[7]_i_6_n_0 ;
  wire \result_reg[8]_i_4_n_0 ;
  wire \result_reg[9]_i_2_n_0 ;
  wire \s_input_ps2_ack[0]_i_1_n_0 ;
  wire \s_input_rs232_rx_ack[0]_i_1_n_0 ;
  wire \s_output_rs232_tx[7]_i_2_n_0 ;
  wire \s_output_rs232_tx[7]_i_3_n_0 ;
  wire \s_output_rs232_tx[7]_i_4_n_0 ;
  wire \s_output_rs232_tx[7]_i_5_n_0 ;
  wire \s_output_rs232_tx[7]_i_6_n_0 ;
  wire \s_output_rs232_tx[7]_i_7_n_0 ;
  wire \s_output_rs232_tx[7]_i_8_n_0 ;
  wire \state[0]_i_1_n_0 ;
  wire \state[1]_i_1_n_0 ;
  wire \state[2]_i_10_n_0 ;
  wire \state[2]_i_11_n_0 ;
  wire \state[2]_i_12_n_0 ;
  wire \state[2]_i_13_n_0 ;
  wire \state[2]_i_14_n_0 ;
  wire \state[2]_i_15_n_0 ;
  wire \state[2]_i_16_n_0 ;
  wire \state[2]_i_17_n_0 ;
  wire \state[2]_i_1_n_0 ;
  wire \state[2]_i_2_n_0 ;
  wire \state[2]_i_3_n_0 ;
  wire \state[2]_i_4_n_0 ;
  wire \state[2]_i_5_n_0 ;
  wire \state[2]_i_6_n_0 ;
  wire \state[2]_i_7_n_0 ;
  wire \state[2]_i_8_n_0 ;
  wire \state[2]_i_9_n_0 ;
  wire \state_reg_n_0_[0] ;
  wire \state_reg_n_0_[1] ;
  wire \state_reg_n_0_[2] ;
  wire [31:0]store_data;
  wire write_enable;
  wire [31:0]write_output;
  wire \write_output[0]_i_1_n_0 ;
  wire \write_output[10]_i_1_n_0 ;
  wire \write_output[11]_i_1_n_0 ;
  wire \write_output[12]_i_1_n_0 ;
  wire \write_output[13]_i_1_n_0 ;
  wire \write_output[14]_i_1_n_0 ;
  wire \write_output[15]_i_1_n_0 ;
  wire \write_output[16]_i_1_n_0 ;
  wire \write_output[17]_i_1_n_0 ;
  wire \write_output[18]_i_1_n_0 ;
  wire \write_output[19]_i_1_n_0 ;
  wire \write_output[1]_i_1_n_0 ;
  wire \write_output[20]_i_1_n_0 ;
  wire \write_output[21]_i_1_n_0 ;
  wire \write_output[22]_i_1_n_0 ;
  wire \write_output[23]_i_1_n_0 ;
  wire \write_output[24]_i_1_n_0 ;
  wire \write_output[25]_i_1_n_0 ;
  wire \write_output[26]_i_1_n_0 ;
  wire \write_output[27]_i_1_n_0 ;
  wire \write_output[28]_i_1_n_0 ;
  wire \write_output[29]_i_1_n_0 ;
  wire \write_output[2]_i_1_n_0 ;
  wire \write_output[30]_i_1_n_0 ;
  wire \write_output[31]_i_1_n_0 ;
  wire \write_output[31]_i_2_n_0 ;
  wire \write_output[31]_i_3_n_0 ;
  wire \write_output[31]_i_4_n_0 ;
  wire \write_output[3]_i_1_n_0 ;
  wire \write_output[4]_i_1_n_0 ;
  wire \write_output[5]_i_1_n_0 ;
  wire \write_output[6]_i_1_n_0 ;
  wire \write_output[7]_i_1_n_0 ;
  wire \write_output[8]_i_1_n_0 ;
  wire \write_output[9]_i_1_n_0 ;
  wire [7:0]write_value;
  wire \write_value[7]_i_3_n_0 ;
  wire NLW_memory_reg_0_CASCADEOUTA_UNCONNECTED;
  wire NLW_memory_reg_0_CASCADEOUTB_UNCONNECTED;
  wire NLW_memory_reg_0_DBITERR_UNCONNECTED;
  wire NLW_memory_reg_0_INJECTDBITERR_UNCONNECTED;
  wire NLW_memory_reg_0_INJECTSBITERR_UNCONNECTED;
  wire NLW_memory_reg_0_REGCEAREGCE_UNCONNECTED;
  wire NLW_memory_reg_0_REGCEB_UNCONNECTED;
  wire NLW_memory_reg_0_SBITERR_UNCONNECTED;
  wire [31:4]NLW_memory_reg_0_DOADO_UNCONNECTED;
  wire [31:0]NLW_memory_reg_0_DOBDO_UNCONNECTED;
  wire [3:0]NLW_memory_reg_0_DOPADOP_UNCONNECTED;
  wire [3:0]NLW_memory_reg_0_DOPBDOP_UNCONNECTED;
  wire [7:0]NLW_memory_reg_0_ECCPARITY_UNCONNECTED;
  wire [8:0]NLW_memory_reg_0_RDADDRECC_UNCONNECTED;
  wire NLW_memory_reg_1_CASCADEOUTA_UNCONNECTED;
  wire NLW_memory_reg_1_CASCADEOUTB_UNCONNECTED;
  wire NLW_memory_reg_1_DBITERR_UNCONNECTED;
  wire NLW_memory_reg_1_INJECTDBITERR_UNCONNECTED;
  wire NLW_memory_reg_1_INJECTSBITERR_UNCONNECTED;
  wire NLW_memory_reg_1_REGCEAREGCE_UNCONNECTED;
  wire NLW_memory_reg_1_REGCEB_UNCONNECTED;
  wire NLW_memory_reg_1_SBITERR_UNCONNECTED;
  wire [31:4]NLW_memory_reg_1_DOADO_UNCONNECTED;
  wire [31:0]NLW_memory_reg_1_DOBDO_UNCONNECTED;
  wire [3:0]NLW_memory_reg_1_DOPADOP_UNCONNECTED;
  wire [3:0]NLW_memory_reg_1_DOPBDOP_UNCONNECTED;
  wire [7:0]NLW_memory_reg_1_ECCPARITY_UNCONNECTED;
  wire [8:0]NLW_memory_reg_1_RDADDRECC_UNCONNECTED;
  wire NLW_memory_reg_2_CASCADEOUTA_UNCONNECTED;
  wire NLW_memory_reg_2_CASCADEOUTB_UNCONNECTED;
  wire NLW_memory_reg_2_DBITERR_UNCONNECTED;
  wire NLW_memory_reg_2_INJECTDBITERR_UNCONNECTED;
  wire NLW_memory_reg_2_INJECTSBITERR_UNCONNECTED;
  wire NLW_memory_reg_2_REGCEAREGCE_UNCONNECTED;
  wire NLW_memory_reg_2_REGCEB_UNCONNECTED;
  wire NLW_memory_reg_2_SBITERR_UNCONNECTED;
  wire [31:4]NLW_memory_reg_2_DOADO_UNCONNECTED;
  wire [31:0]NLW_memory_reg_2_DOBDO_UNCONNECTED;
  wire [3:0]NLW_memory_reg_2_DOPADOP_UNCONNECTED;
  wire [3:0]NLW_memory_reg_2_DOPBDOP_UNCONNECTED;
  wire [7:0]NLW_memory_reg_2_ECCPARITY_UNCONNECTED;
  wire [8:0]NLW_memory_reg_2_RDADDRECC_UNCONNECTED;
  wire NLW_memory_reg_3_CASCADEOUTA_UNCONNECTED;
  wire NLW_memory_reg_3_CASCADEOUTB_UNCONNECTED;
  wire NLW_memory_reg_3_DBITERR_UNCONNECTED;
  wire NLW_memory_reg_3_INJECTDBITERR_UNCONNECTED;
  wire NLW_memory_reg_3_INJECTSBITERR_UNCONNECTED;
  wire NLW_memory_reg_3_REGCEAREGCE_UNCONNECTED;
  wire NLW_memory_reg_3_REGCEB_UNCONNECTED;
  wire NLW_memory_reg_3_SBITERR_UNCONNECTED;
  wire [31:4]NLW_memory_reg_3_DOADO_UNCONNECTED;
  wire [31:0]NLW_memory_reg_3_DOBDO_UNCONNECTED;
  wire [3:0]NLW_memory_reg_3_DOPADOP_UNCONNECTED;
  wire [3:0]NLW_memory_reg_3_DOPBDOP_UNCONNECTED;
  wire [7:0]NLW_memory_reg_3_ECCPARITY_UNCONNECTED;
  wire [8:0]NLW_memory_reg_3_RDADDRECC_UNCONNECTED;
  wire NLW_memory_reg_4_CASCADEOUTA_UNCONNECTED;
  wire NLW_memory_reg_4_CASCADEOUTB_UNCONNECTED;
  wire NLW_memory_reg_4_DBITERR_UNCONNECTED;
  wire NLW_memory_reg_4_INJECTDBITERR_UNCONNECTED;
  wire NLW_memory_reg_4_INJECTSBITERR_UNCONNECTED;
  wire NLW_memory_reg_4_REGCEAREGCE_UNCONNECTED;
  wire NLW_memory_reg_4_REGCEB_UNCONNECTED;
  wire NLW_memory_reg_4_SBITERR_UNCONNECTED;
  wire [31:4]NLW_memory_reg_4_DOADO_UNCONNECTED;
  wire [31:0]NLW_memory_reg_4_DOBDO_UNCONNECTED;
  wire [3:0]NLW_memory_reg_4_DOPADOP_UNCONNECTED;
  wire [3:0]NLW_memory_reg_4_DOPBDOP_UNCONNECTED;
  wire [7:0]NLW_memory_reg_4_ECCPARITY_UNCONNECTED;
  wire [8:0]NLW_memory_reg_4_RDADDRECC_UNCONNECTED;
  wire NLW_memory_reg_5_CASCADEOUTA_UNCONNECTED;
  wire NLW_memory_reg_5_CASCADEOUTB_UNCONNECTED;
  wire NLW_memory_reg_5_DBITERR_UNCONNECTED;
  wire NLW_memory_reg_5_INJECTDBITERR_UNCONNECTED;
  wire NLW_memory_reg_5_INJECTSBITERR_UNCONNECTED;
  wire NLW_memory_reg_5_REGCEAREGCE_UNCONNECTED;
  wire NLW_memory_reg_5_REGCEB_UNCONNECTED;
  wire NLW_memory_reg_5_SBITERR_UNCONNECTED;
  wire [31:4]NLW_memory_reg_5_DOADO_UNCONNECTED;
  wire [31:0]NLW_memory_reg_5_DOBDO_UNCONNECTED;
  wire [3:0]NLW_memory_reg_5_DOPADOP_UNCONNECTED;
  wire [3:0]NLW_memory_reg_5_DOPBDOP_UNCONNECTED;
  wire [7:0]NLW_memory_reg_5_ECCPARITY_UNCONNECTED;
  wire [8:0]NLW_memory_reg_5_RDADDRECC_UNCONNECTED;
  wire NLW_memory_reg_6_CASCADEOUTA_UNCONNECTED;
  wire NLW_memory_reg_6_CASCADEOUTB_UNCONNECTED;
  wire NLW_memory_reg_6_DBITERR_UNCONNECTED;
  wire NLW_memory_reg_6_INJECTDBITERR_UNCONNECTED;
  wire NLW_memory_reg_6_INJECTSBITERR_UNCONNECTED;
  wire NLW_memory_reg_6_REGCEAREGCE_UNCONNECTED;
  wire NLW_memory_reg_6_REGCEB_UNCONNECTED;
  wire NLW_memory_reg_6_SBITERR_UNCONNECTED;
  wire [31:4]NLW_memory_reg_6_DOADO_UNCONNECTED;
  wire [31:0]NLW_memory_reg_6_DOBDO_UNCONNECTED;
  wire [3:0]NLW_memory_reg_6_DOPADOP_UNCONNECTED;
  wire [3:0]NLW_memory_reg_6_DOPBDOP_UNCONNECTED;
  wire [7:0]NLW_memory_reg_6_ECCPARITY_UNCONNECTED;
  wire [8:0]NLW_memory_reg_6_RDADDRECC_UNCONNECTED;
  wire NLW_memory_reg_7_CASCADEOUTA_UNCONNECTED;
  wire NLW_memory_reg_7_CASCADEOUTB_UNCONNECTED;
  wire NLW_memory_reg_7_DBITERR_UNCONNECTED;
  wire NLW_memory_reg_7_INJECTDBITERR_UNCONNECTED;
  wire NLW_memory_reg_7_INJECTSBITERR_UNCONNECTED;
  wire NLW_memory_reg_7_REGCEAREGCE_UNCONNECTED;
  wire NLW_memory_reg_7_REGCEB_UNCONNECTED;
  wire NLW_memory_reg_7_SBITERR_UNCONNECTED;
  wire [31:4]NLW_memory_reg_7_DOADO_UNCONNECTED;
  wire [31:0]NLW_memory_reg_7_DOBDO_UNCONNECTED;
  wire [3:0]NLW_memory_reg_7_DOPADOP_UNCONNECTED;
  wire [3:0]NLW_memory_reg_7_DOPBDOP_UNCONNECTED;
  wire [7:0]NLW_memory_reg_7_ECCPARITY_UNCONNECTED;
  wire [8:0]NLW_memory_reg_7_RDADDRECC_UNCONNECTED;
  wire [3:0]\NLW_program_counter_reg[15]_i_3_CO_UNCONNECTED ;
  wire [3:3]\NLW_program_counter_reg[15]_i_3_O_UNCONNECTED ;
  wire [2:0]\NLW_program_counter_reg_rep[4]_i_2_CO_UNCONNECTED ;
  wire [2:0]\NLW_program_counter_reg_rep[8]_i_2_CO_UNCONNECTED ;
  wire [2:0]\NLW_program_counter_reg_rep[9]_i_5_CO_UNCONNECTED ;
  wire [1:0]NLW_registers_reg_r1_0_15_0_5_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r1_0_15_12_17_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r1_0_15_18_23_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r1_0_15_24_29_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r1_0_15_30_31_DOB_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r1_0_15_30_31_DOC_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r1_0_15_30_31_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r1_0_15_6_11_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r2_0_15_0_5_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r2_0_15_12_17_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r2_0_15_18_23_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r2_0_15_24_29_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r2_0_15_30_31_DOB_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r2_0_15_30_31_DOC_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r2_0_15_30_31_DOD_UNCONNECTED;
  wire [1:0]NLW_registers_reg_r2_0_15_6_11_DOD_UNCONNECTED;
  wire [2:0]\NLW_result_reg[0]_i_11_CO_UNCONNECTED ;
  wire [3:0]\NLW_result_reg[0]_i_11_O_UNCONNECTED ;
  wire [3:0]\NLW_result_reg[0]_i_4_CO_UNCONNECTED ;
  wire [3:0]\NLW_result_reg[0]_i_4_O_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[0]_i_7_CO_UNCONNECTED ;
  wire [3:0]\NLW_result_reg[0]_i_7_O_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[11]_i_4_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[11]_i_5_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[11]_i_6_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[12]_i_3_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[15]_i_2_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[16]_i_4_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[16]_i_6_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[16]_i_8_CO_UNCONNECTED ;
  wire [3:3]\NLW_result_reg[16]_i_8_O_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[16]_i_9_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[19]_i_2_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[19]_i_4_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[23]_i_2_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[23]_i_8_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[23]_i_9_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[27]_i_2_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[27]_i_8_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[27]_i_9_CO_UNCONNECTED ;
  wire [3:0]\NLW_result_reg[31]_i_16_CO_UNCONNECTED ;
  wire [3:0]\NLW_result_reg[31]_i_17_CO_UNCONNECTED ;
  wire [3:0]\NLW_result_reg[31]_i_8_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[3]_i_3_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[3]_i_5_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[3]_i_6_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[4]_i_4_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[7]_i_3_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[7]_i_6_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[8]_i_4_CO_UNCONNECTED ;
  wire [2:0]\NLW_result_reg[9]_i_2_CO_UNCONNECTED ;
  FDRE \address_a_2_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(address_a[0]),
        .Q(address_a_2[0]),
        .R(1'b0));
  FDRE \address_a_2_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(address_a[1]),
        .Q(address_a_2[1]),
        .R(1'b0));
  FDRE \address_a_2_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(address_a[2]),
        .Q(address_a_2[2]),
        .R(1'b0));
  FDRE \address_a_2_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(address_a[3]),
        .Q(address_a_2[3]),
        .R(1'b0));
  FDRE \address_b_2_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[0] ),
        .Q(address_b_2[0]),
        .R(1'b0));
  FDRE \address_b_2_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[1] ),
        .Q(address_b_2[1]),
        .R(1'b0));
  FDRE \address_b_2_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[2] ),
        .Q(address_b_2[2]),
        .R(1'b0));
  FDRE \address_b_2_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[3] ),
        .Q(address_b_2[3]),
        .R(1'b0));
  FDRE \address_z_2_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(address_z[0]),
        .Q(address_z_2[0]),
        .R(1'b0));
  FDRE \address_z_2_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(address_z[1]),
        .Q(address_z_2[1]),
        .R(1'b0));
  FDRE \address_z_2_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(address_z[2]),
        .Q(address_z_2[2]),
        .R(1'b0));
  FDRE \address_z_2_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(address_z[3]),
        .Q(address_z_2[3]),
        .R(1'b0));
  LUT3 #(
    .INIT(8'h20))
    \address_z_3[3]_i_1
       (.I0(\state_reg_n_0_[0] ),
        .I1(\state_reg_n_0_[2] ),
        .I2(\state_reg_n_0_[1] ),
        .O(\address_z_3[3]_i_1_n_0 ));
  FDRE \address_z_3_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(\address_z_3[3]_i_1_n_0 ),
        .D(address_z_2[0]),
        .Q(address_z_3[0]),
        .R(INTERNAL_RST_reg));
  FDRE \address_z_3_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(\address_z_3[3]_i_1_n_0 ),
        .D(address_z_2[1]),
        .Q(address_z_3[1]),
        .R(INTERNAL_RST_reg));
  FDRE \address_z_3_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(\address_z_3[3]_i_1_n_0 ),
        .D(address_z_2[2]),
        .Q(address_z_3[2]),
        .R(INTERNAL_RST_reg));
  FDRE \address_z_3_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(\address_z_3[3]_i_1_n_0 ),
        .D(address_z_2[3]),
        .Q(address_z_3[3]),
        .R(INTERNAL_RST_reg));
  LUT6 #(
    .INIT(64'hFFDF55DFFFDFFFDF))
    \instruction[0]_i_1
       (.I0(\instruction_reg[0]_i_2_n_0 ),
        .I1(\instruction[0]_i_3_n_0 ),
        .I2(\instruction_reg[0]_i_4_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction_reg[0]_i_5_n_0 ),
        .I5(\instruction[0]_i_6_n_0 ),
        .O(\instruction[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004F40404))
    \instruction[0]_i_11
       (.I0(\instruction_reg[0]_i_24_n_0 ),
        .I1(\instruction[0]_i_25_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\instruction[0]_i_26_n_0 ),
        .I4(\instruction_reg[0]_i_27_n_0 ),
        .I5(\instruction[0]_i_28_n_0 ),
        .O(\instruction[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8A8AA8AAA8AAA8AA))
    \instruction[0]_i_12
       (.I0(\instruction[0]_i_29_n_0 ),
        .I1(\instruction[0]_i_30_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[0]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAA800008))
    \instruction[0]_i_13
       (.I0(\instruction[0]_i_31_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00040004FFFF0000))
    \instruction[0]_i_14
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\instruction[7]_i_17_n_0 ),
        .I4(\instruction[0]_i_32_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[0]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h00002EEE))
    \instruction[0]_i_15
       (.I0(\instruction_reg[0]_i_33_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[0]_i_34_n_0 ),
        .I3(\instruction[0]_i_35_n_0 ),
        .I4(\instruction_reg[0]_i_36_n_0 ),
        .O(\instruction[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA02F20AFA02020))
    \instruction[0]_i_16
       (.I0(\instruction_reg[0]_i_37_n_0 ),
        .I1(\instruction[0]_i_38_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\instruction_reg[0]_i_39_n_0 ),
        .I4(\instruction[7]_i_17_n_0 ),
        .I5(\instruction[0]_i_40_n_0 ),
        .O(\instruction[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hC000003038000804))
    \instruction[0]_i_17
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBDEEFF7DFFFFFFFF))
    \instruction[0]_i_18
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[0]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h08000214))
    \instruction[0]_i_19
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[0]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h00240000))
    \instruction[0]_i_21
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000800))
    \instruction[0]_i_22
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h1A00004000000040))
    \instruction[0]_i_23
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFFFEFFFF))
    \instruction[0]_i_25
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0002A0800A140000))
    \instruction[0]_i_26
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000300044000000))
    \instruction[0]_i_28
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\instruction[26]_i_17_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hA800A800A8FFA800))
    \instruction[0]_i_29
       (.I0(\instruction_reg[0]_i_47_n_0 ),
        .I1(\instruction[25]_i_15_n_0 ),
        .I2(\instruction[0]_i_48_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\instruction[0]_i_49_n_0 ),
        .I5(\instruction_reg[0]_i_50_n_0 ),
        .O(\instruction[0]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h28FF2800))
    \instruction[0]_i_3
       (.I0(\instruction[0]_i_9_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\instruction_reg[0]_i_10_n_0 ),
        .O(\instruction[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEFFFFFFFFFFAB))
    \instruction[0]_i_30
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[0]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'h0A004520))
    \instruction[0]_i_31
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004042110))
    \instruction[0]_i_32
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[0]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h00F000400F00F00F))
    \instruction[0]_i_34
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAEAAFF))
    \instruction[0]_i_35
       (.I0(\instruction[0]_i_53_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\instruction[0]_i_48_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[0]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h08))
    \instruction[0]_i_38
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hF7))
    \instruction[0]_i_40
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[0]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDFFD575FFF7F))
    \instruction[0]_i_41
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFADFFFFFFFFFFF))
    \instruction[0]_i_42
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h3030030C3CA8C088))
    \instruction[0]_i_43
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[0]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h000000004A042944))
    \instruction[0]_i_44
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[0]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h7F7FBCA97F7FBFEB))
    \instruction[0]_i_45
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[0]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hE4F5BEAAEEFFB6F7))
    \instruction[0]_i_46
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[0]_i_46_n_0 ));
  LUT3 #(
    .INIT(8'hFB))
    \instruction[0]_i_48
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[0]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h7F7F3FFFFFFFFFF7))
    \instruction[0]_i_49
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDFFDDFFFDF2DD))
    \instruction[0]_i_51
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[0]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEFEFFFFEFFEFF))
    \instruction[0]_i_52
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[0]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000))
    \instruction[0]_i_53
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[0]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0000040404000000))
    \instruction[0]_i_54
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000898100))
    \instruction[0]_i_55
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[0]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFCFFFCBBFB))
    \instruction[0]_i_56
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[0]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h7F007F7F7FBF7FBF))
    \instruction[0]_i_57
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFFFFFFEFFEFF))
    \instruction[0]_i_58
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[0]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7F7FBBFC7FBB))
    \instruction[0]_i_59
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[0]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888B8B8B8B8))
    \instruction[0]_i_6
       (.I0(\instruction[0]_i_15_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\instruction[0]_i_16_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\instruction[6]_i_13_n_0 ),
        .I5(\instruction[0]_i_17_n_0 ),
        .O(\instruction[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFEDFFB7EFFFEFEF))
    \instruction[0]_i_60
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[0]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFFCFEF3EEEF033CF))
    \instruction[0]_i_61
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[0]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h2248214A41004091))
    \instruction[0]_i_62
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[0]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h00AAA50025100210))
    \instruction[0]_i_63
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[0]_i_63_n_0 ));
  LUT5 #(
    .INIT(32'hBB8BBBBB))
    \instruction[0]_i_7
       (.I0(\instruction[0]_i_18_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\instruction[0]_i_19_n_0 ),
        .O(\instruction[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h8B8BBBBBBBBBBB8B))
    \instruction[0]_i_8
       (.I0(\instruction_reg[0]_i_20_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[0]_i_21_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h02495A0000200002))
    \instruction[0]_i_9
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hBB8B8888BB8BBBBB))
    \instruction[15]_i_1
       (.I0(\instruction[15]_i_2_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[15]_i_3_n_0 ),
        .I3(\instruction[15]_i_4_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction[15]_i_5_n_0 ),
        .O(\instruction[15]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h4E444454))
    \instruction[15]_i_10
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF))
    \instruction[15]_i_11
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h3FF7FBFB3FFFFFFF))
    \instruction[15]_i_12
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hEE44444481100010))
    \instruction[15]_i_13
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF))
    \instruction[15]_i_14
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep_n_0_[0] ),
        .O(\instruction[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF1FFFFF7F7FFF))
    \instruction[15]_i_15
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[15]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFF5FFFFEEFBFFFF))
    \instruction[15]_i_16
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[15]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFFFFFFFF3F7FFF7))
    \instruction[15]_i_17
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[15]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h4010401F))
    \instruction[15]_i_18
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8880FFFF88800000))
    \instruction[15]_i_2
       (.I0(\instruction[15]_i_6_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\instruction[15]_i_7_n_0 ),
        .O(\instruction[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBB8BBBBBBBBBB))
    \instruction[15]_i_3
       (.I0(\instruction[15]_i_8_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\instruction[15]_i_9_n_0 ),
        .I5(\instruction[15]_i_10_n_0 ),
        .O(\instruction[15]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h8000))
    \instruction[15]_i_4
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB800B8FFB8FFB8FF))
    \instruction[15]_i_5
       (.I0(\instruction[15]_i_11_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\instruction[15]_i_12_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\instruction[15]_i_13_n_0 ),
        .O(\instruction[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4000004108020041))
    \instruction[15]_i_6
       (.I0(\program_counter_reg_rep_n_0_[0] ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h575757F7F7F757F7))
    \instruction[15]_i_7
       (.I0(\instruction[15]_i_14_n_0 ),
        .I1(\instruction[15]_i_15_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\instruction[15]_i_16_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction[15]_i_17_n_0 ),
        .O(\instruction[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h07FFFFFF))
    \instruction[15]_i_8
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\instruction[15]_i_18_n_0 ),
        .O(\instruction[15]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[15]_i_9
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00EAFFEAFFFFFFFF))
    \instruction[16]_i_1
       (.I0(\instruction[16]_i_2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\instruction_reg[16]_i_3_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\instruction[16]_i_4_n_0 ),
        .I5(\instruction_reg[16]_i_5_n_0 ),
        .O(\instruction[16]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hD5DDFFFFD5DD0000))
    \instruction[16]_i_10
       (.I0(\instruction[16]_i_14_n_0 ),
        .I1(\instruction[16]_i_15_n_0 ),
        .I2(\instruction[16]_i_16_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\instruction_reg[16]_i_17_n_0 ),
        .O(\instruction[16]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[16]_i_11
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[16]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00002A00))
    \instruction[16]_i_12
       (.I0(\instruction_reg[16]_i_18_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\instruction[16]_i_19_n_0 ),
        .I3(\instruction[16]_i_20_n_0 ),
        .I4(\instruction[16]_i_21_n_0 ),
        .O(\instruction[16]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000000000A8A2AAA))
    \instruction[16]_i_13
       (.I0(\instruction_reg[16]_i_22_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\instruction[16]_i_23_n_0 ),
        .I4(\instruction[16]_i_24_n_0 ),
        .I5(\instruction[16]_i_25_n_0 ),
        .O(\instruction[16]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE))
    \instruction[16]_i_14
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFEEFFEEE5))
    \instruction[16]_i_15
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h7F))
    \instruction[16]_i_16
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[16]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h002880E004200040))
    \instruction[16]_i_19
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF0400000404))
    \instruction[16]_i_2
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\instruction[16]_i_6_n_0 ),
        .I3(\instruction[16]_i_7_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[1] ),
        .O(\instruction[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFCFDDFFFF))
    \instruction[16]_i_20
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\instruction[7]_i_12_n_0 ),
        .O(\instruction[16]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h202022220000FF00))
    \instruction[16]_i_21
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\instruction[7]_i_12_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\instruction[16]_i_7_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[16]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h3C08000000008080))
    \instruction[16]_i_23
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h00800280))
    \instruction[16]_i_24
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080))
    \instruction[16]_i_25
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[16]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFFFFFFFFFDFFD))
    \instruction[16]_i_26
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[16]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFD5D5DFDFFFF7FFF))
    \instruction[16]_i_27
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[16]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hBBBB8BBBBBBBBBBB))
    \instruction[16]_i_28
       (.I0(\instruction[16]_i_32_n_0 ),
        .I1(\instruction[16]_i_33_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[16]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFF700F7))
    \instruction[16]_i_29
       (.I0(\instruction[16]_i_34_n_0 ),
        .I1(\instruction[16]_i_35_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\instruction[16]_i_36_n_0 ),
        .I5(\instruction[16]_i_37_n_0 ),
        .O(\instruction[16]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010501F5F))
    \instruction[16]_i_30
       (.I0(\instruction[16]_i_38_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\instruction[16]_i_39_n_0 ),
        .I4(\instruction[16]_i_40_n_0 ),
        .I5(\instruction[16]_i_37_n_0 ),
        .O(\instruction[16]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h5DDDDDDD5DDD5555))
    \instruction[16]_i_31
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\instruction[16]_i_41_n_0 ),
        .I2(\instruction[21]_i_30_n_0 ),
        .I3(\instruction[16]_i_34_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\instruction[16]_i_42_n_0 ),
        .O(\instruction[16]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFF9867FF))
    \instruction[16]_i_32
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h85800D0000002E40))
    \instruction[16]_i_33
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[16]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h01))
    \instruction[16]_i_34
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[16]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h01))
    \instruction[16]_i_35
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h7CFF7C00))
    \instruction[16]_i_36
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\instruction[16]_i_43_n_0 ),
        .I4(\instruction[16]_i_44_n_0 ),
        .O(\instruction[16]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000))
    \instruction[16]_i_37
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[16]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0000880000411110))
    \instruction[16]_i_38
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[16]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h00083374))
    \instruction[16]_i_39
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[16]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA8AAAAAA))
    \instruction[16]_i_4
       (.I0(\instruction[16]_i_10_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\instruction[16]_i_11_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000))
    \instruction[16]_i_40
       (.I0(\instruction[16]_i_45_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFF72BFFF))
    \instruction[16]_i_41
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[16]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h00FFFFDFFFFF8F8F))
    \instruction[16]_i_42
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[16]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'h04040914))
    \instruction[16]_i_43
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[16]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h00D7F7D7D7F7D7F7))
    \instruction[16]_i_44
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[2] ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[16]_i_44_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[16]_i_45
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[16]_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[16]_i_6
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[16]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h8000))
    \instruction[16]_i_7
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0054A01A0150000A))
    \instruction[16]_i_8
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h000F000040104010))
    \instruction[16]_i_9
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[16]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF5F555D5FFFFFFFF))
    \instruction[17]_i_1
       (.I0(\instruction[17]_i_2_n_0 ),
        .I1(\instruction_reg[17]_i_3_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\instruction_reg[17]_i_4_n_0 ),
        .I5(\instruction[17]_i_5_n_0 ),
        .O(\instruction[17]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h3200F00101C00200))
    \instruction[17]_i_10
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[17]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hA004AA1210200098))
    \instruction[17]_i_11
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[17]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00A1FFFF00A10000))
    \instruction[17]_i_13
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\instruction[17]_i_19_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\instruction[17]_i_20_n_0 ),
        .O(\instruction[17]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h44FC74FC74FC74FC))
    \instruction[17]_i_15
       (.I0(\instruction[17]_i_23_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[17]_i_24_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\instruction[17]_i_25_n_0 ),
        .O(\instruction[17]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7FFFFFF))
    \instruction[17]_i_16
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[17]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000A0A2A8AA))
    \instruction[17]_i_17
       (.I0(\instruction_reg[17]_i_26_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\instruction[17]_i_27_n_0 ),
        .I4(\instruction[17]_i_28_n_0 ),
        .I5(\instruction[17]_i_29_n_0 ),
        .O(\instruction[17]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022E2EEE2))
    \instruction[17]_i_18
       (.I0(\instruction_reg[17]_i_30_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[17]_i_31_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\instruction[17]_i_32_n_0 ),
        .I5(\instruction[17]_i_33_n_0 ),
        .O(\instruction[17]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hE6E6E6FFFFFFFFFF))
    \instruction[17]_i_19
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[17]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFFFFF00FFFFFF))
    \instruction[17]_i_2
       (.I0(\instruction[17]_i_6_n_0 ),
        .I1(\instruction[17]_i_7_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\instruction[25]_i_7_n_0 ),
        .O(\instruction[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000024000000))
    \instruction[17]_i_20
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\instruction[23]_i_22_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[17]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEE222E2))
    \instruction[17]_i_21
       (.I0(\instruction[17]_i_34_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[17]_i_31_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\instruction[17]_i_35_n_0 ),
        .I5(\instruction[17]_i_36_n_0 ),
        .O(\instruction[17]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2))
    \instruction[17]_i_22
       (.I0(\instruction[17]_i_37_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\instruction[17]_i_38_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\instruction[17]_i_39_n_0 ),
        .I5(\instruction[17]_i_40_n_0 ),
        .O(\instruction[17]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h48FF6AEE48006A22))
    \instruction[17]_i_23
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[17]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBB8))
    \instruction[17]_i_24
       (.I0(\instruction[17]_i_41_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\instruction[7]_i_12_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[17]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h24))
    \instruction[17]_i_25
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[17]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000028424014))
    \instruction[17]_i_27
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[17]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h000101000000D020))
    \instruction[17]_i_28
       (.I0(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[17]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h8080000000008088))
    \instruction[17]_i_29
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[17]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFBBEEFFBBEEF))
    \instruction[17]_i_31
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[17]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hD6018141D6018168))
    \instruction[17]_i_32
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[17]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0380000))
    \instruction[17]_i_33
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\instruction[23]_i_22_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[17]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA2AAAAAAA))
    \instruction[17]_i_34
       (.I0(\instruction_reg[17]_i_46_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[17]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hCCBFCBFCFFCBFCBF))
    \instruction[17]_i_35
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[17]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0800000000000400))
    \instruction[17]_i_36
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\instruction[23]_i_22_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[17]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hDFF5DAEFDAEFF5DA))
    \instruction[17]_i_37
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[17]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFADADFAFADFFFED))
    \instruction[17]_i_38
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[17]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBAB888888A8))
    \instruction[17]_i_39
       (.I0(\instruction[17]_i_47_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\instruction[17]_i_48_n_0 ),
        .I5(\instruction[17]_i_49_n_0 ),
        .O(\instruction[17]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0440000400000000))
    \instruction[17]_i_40
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\instruction[23]_i_22_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[17]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h477F0FF7FFFFFEFF))
    \instruction[17]_i_41
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[17]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h56DB6DB6FFEDFFFF))
    \instruction[17]_i_42
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[17]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h9B9E9FF7EF7D5D9E))
    \instruction[17]_i_43
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[17]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hEEFDEFDEF5EFDEFD))
    \instruction[17]_i_44
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[17]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hBBFDFD46F6BBB95D))
    \instruction[17]_i_45
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[17]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hEFDE5567FEFF6756))
    \instruction[17]_i_47
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[17]_i_47_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[17]_i_48
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[17]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFFB79BE9ECFE7))
    \instruction[17]_i_49
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[17]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h2F20202020202020))
    \instruction[17]_i_5
       (.I0(\instruction_reg[17]_i_12_n_0 ),
        .I1(\instruction[17]_i_13_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[0] ),
        .I3(\instruction_reg[17]_i_14_n_0 ),
        .I4(\instruction[17]_i_15_n_0 ),
        .I5(\instruction[17]_i_16_n_0 ),
        .O(\instruction[17]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hECE31FDC2FFEEB3F))
    \instruction[17]_i_50
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[17]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFBFEFFEBFEBFABFE))
    \instruction[17]_i_51
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[17]_i_51_n_0 ));
  LUT5 #(
    .INIT(32'h44083330))
    \instruction[17]_i_6
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[17]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[17]_i_7
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4010020048180110))
    \instruction[17]_i_8
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h24765A806426008D))
    \instruction[17]_i_9
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[17]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h575757F7F7F757F7))
    \instruction[18]_i_1
       (.I0(\instruction[18]_i_2_n_0 ),
        .I1(\instruction[18]_i_3_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\instruction_reg[18]_i_4_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction_reg[18]_i_5_n_0 ),
        .O(\instruction[18]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F4040000))
    \instruction[18]_i_11
       (.I0(\instruction[18]_i_24_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[2] ),
        .I3(\instruction[18]_i_25_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I5(\instruction[18]_i_26_n_0 ),
        .O(\instruction[18]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF4F70407F4F7F4F7))
    \instruction[18]_i_14
       (.I0(\instruction[18]_i_31_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\instruction[18]_i_32_n_0 ),
        .I3(\instruction[18]_i_33_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\instruction[18]_i_34_n_0 ),
        .O(\instruction[18]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00E2E2E2E2E2E2E2))
    \instruction[18]_i_15
       (.I0(\instruction[18]_i_35_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\instruction[18]_i_36_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[18]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h2816148000000000))
    \instruction[18]_i_16
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0224408202900000))
    \instruction[18]_i_17
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h000057F7FFFF57F7))
    \instruction[18]_i_18
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[18]_i_19
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[18]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFBBBFBFBFBF))
    \instruction[18]_i_2
       (.I0(\instruction[18]_i_6_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction[18]_i_7_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFAAFFEFF))
    \instruction[18]_i_20
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[18]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h07))
    \instruction[18]_i_24
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h0020))
    \instruction[18]_i_25
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[18]_i_26
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[18]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h7275EBFF7567DE7F))
    \instruction[18]_i_27
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[18]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFEED5FFEDF7FEDFF))
    \instruction[18]_i_28
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFF19B95EFEF7EFEF))
    \instruction[18]_i_29
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h0000F404))
    \instruction[18]_i_3
       (.I0(\instruction_reg[18]_i_8_n_0 ),
        .I1(\instruction[18]_i_9_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[0] ),
        .I3(\instruction_reg[18]_i_10_n_0 ),
        .I4(\instruction[18]_i_11_n_0 ),
        .O(\instruction[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h675E75FF75EF56FF))
    \instruction[18]_i_30
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[18]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'h18846018))
    \instruction[18]_i_31
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[18]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h8A))
    \instruction[18]_i_32
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h01486804))
    \instruction[18]_i_33
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[18]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'h0010))
    \instruction[18]_i_34
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[18]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFEBFBFEFFFEBEFFF))
    \instruction[18]_i_35
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[18]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFEFDEFD7F5E75EF7))
    \instruction[18]_i_36
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[18]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF6D6BDFFFF))
    \instruction[18]_i_37
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFBEBEF7F77FFB7F))
    \instruction[18]_i_38
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[18]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hBBBDD66BD6FFBDFF))
    \instruction[18]_i_39
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[18]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hEEEFEFEFFFFFFFFE))
    \instruction[18]_i_40
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[18]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFEFBFBEFEFBEF75F))
    \instruction[18]_i_41
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFEE55FFEDFFFE5FF))
    \instruction[18]_i_42
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[18]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[18]_i_6
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[18]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[18]_i_7
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFB08FFFFFB080000))
    \instruction[18]_i_9
       (.I0(\instruction[18]_i_18_n_0 ),
        .I1(\instruction[18]_i_19_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[2] ),
        .I3(\instruction[18]_i_20_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\instruction_reg[18]_i_21_n_0 ),
        .O(\instruction[18]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFF8F888FFF8FFF8F))
    \instruction[19]_i_1
       (.I0(\instruction[19]_i_2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\instruction[19]_i_3_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction[19]_i_4_n_0 ),
        .I5(\instruction[19]_i_5_n_0 ),
        .O(\instruction[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h40000000))
    \instruction[19]_i_11
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[19]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hDDFFFFFD))
    \instruction[19]_i_13
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[19]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h7777777747777777))
    \instruction[19]_i_14
       (.I0(\instruction[19]_i_23_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\instruction[19]_i_24_n_0 ),
        .I4(\instruction[19]_i_25_n_0 ),
        .I5(\instruction[19]_i_26_n_0 ),
        .O(\instruction[19]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBEAEFFFBFBFFF))
    \instruction[19]_i_15
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[19]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFF5ABF7FFFFFFF7))
    \instruction[19]_i_16
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[19]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001A40))
    \instruction[19]_i_17
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[19]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[19]_i_18
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[19]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFE6FF))
    \instruction[19]_i_19
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[19]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hB800B800B8FFB800))
    \instruction[19]_i_2
       (.I0(\instruction[19]_i_6_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[19]_i_7_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\instruction[19]_i_8_n_0 ),
        .O(\instruction[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h7777F77FF3FFFFFF))
    \instruction[19]_i_20
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[19]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h5FFDFDFD))
    \instruction[19]_i_21
       (.I0(\instruction[19]_i_27_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[19]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFF6DFFFF))
    \instruction[19]_i_22
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\instruction[19]_i_28_n_0 ),
        .O(\instruction[19]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h02FFFFFFFFFFFFFF))
    \instruction[19]_i_23
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\instruction[19]_i_29_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\instruction[19]_i_30_n_0 ),
        .I4(\instruction[19]_i_31_n_0 ),
        .I5(\instruction[19]_i_32_n_0 ),
        .O(\instruction[19]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h6))
    \instruction[19]_i_24
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .O(\instruction[19]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[19]_i_25
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[19]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h6))
    \instruction[19]_i_26
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[19]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h30303000888888B8))
    \instruction[19]_i_27
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[19]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h00982200))
    \instruction[19]_i_28
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[19]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h7F))
    \instruction[19]_i_29
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[19]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000))
    \instruction[19]_i_3
       (.I0(\instruction[19]_i_9_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\instruction_reg[19]_i_10_n_0 ),
        .I3(\instruction[19]_i_11_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\instruction_reg[19]_i_12_n_0 ),
        .O(\instruction[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF))
    \instruction[19]_i_30
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[19]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAFAAEFFFFFFFFFFF))
    \instruction[19]_i_31
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\instruction[25]_i_28_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[19]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBFFFEFFEBFFF))
    \instruction[19]_i_32
       (.I0(\instruction[16]_i_11_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[19]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004E200E2))
    \instruction[19]_i_4
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\instruction[19]_i_13_n_0 ),
        .O(\instruction[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h8B8B8B8BBB8B8B8B))
    \instruction[19]_i_5
       (.I0(\instruction[19]_i_14_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\instruction[19]_i_15_n_0 ),
        .I4(\instruction[19]_i_16_n_0 ),
        .I5(\instruction[19]_i_17_n_0 ),
        .O(\instruction[19]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00004000))
    \instruction[19]_i_6
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200000410))
    \instruction[19]_i_7
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDEFEFFFFEFE7F))
    \instruction[19]_i_8
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF77FFFFF7FFFF))
    \instruction[19]_i_9
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\instruction[19]_i_18_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[1] ),
        .O(\instruction[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h111DDD1DFFFFFFFF))
    \instruction[1]_i_1
       (.I0(\instruction_reg[1]_i_2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\instruction[1]_i_3_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\instruction_reg[1]_i_4_n_0 ),
        .I5(\instruction_reg[1]_i_5_n_0 ),
        .O(\instruction[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004F40404))
    \instruction[1]_i_10
       (.I0(\instruction[1]_i_16_n_0 ),
        .I1(\instruction_reg[1]_i_17_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\instruction_reg[1]_i_18_n_0 ),
        .I4(\instruction[1]_i_19_n_0 ),
        .I5(\instruction[1]_i_20_n_0 ),
        .O(\instruction[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004F40404))
    \instruction[1]_i_11
       (.I0(\instruction[1]_i_21_n_0 ),
        .I1(\instruction[1]_i_22_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\instruction_reg[1]_i_23_n_0 ),
        .I4(\instruction_reg[1]_i_24_n_0 ),
        .I5(\instruction[1]_i_25_n_0 ),
        .O(\instruction[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFEFFBFFFFFFBF))
    \instruction[1]_i_12
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFDFFFF))
    \instruction[1]_i_13
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h734FFFFF7F7FFFFF))
    \instruction[1]_i_14
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFFFFFFFE))
    \instruction[1]_i_15
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020040000))
    \instruction[1]_i_16
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\instruction[20]_i_3_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\instruction[1]_i_26_n_0 ),
        .O(\instruction[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8888888888888))
    \instruction[1]_i_19
       (.I0(\instruction[1]_i_31_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[1]_i_32_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\instruction[1]_i_33_n_0 ),
        .I5(\instruction[1]_i_34_n_0 ),
        .O(\instruction[1]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888))
    \instruction[1]_i_20
       (.I0(\instruction[1]_i_35_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[1]_i_36_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\instruction[1]_i_37_n_0 ),
        .O(\instruction[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000))
    \instruction[1]_i_21
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\instruction[3]_i_23_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h88888888BBB888B8))
    \instruction[1]_i_22
       (.I0(\instruction[1]_i_38_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[1]_i_39_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\instruction[1]_i_40_n_0 ),
        .I5(\instruction[1]_i_41_n_0 ),
        .O(\instruction[1]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h7400740074337400))
    \instruction[1]_i_25
       (.I0(\instruction[1]_i_46_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[1]_i_47_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\instruction[24]_i_27_n_0 ),
        .I5(\instruction[7]_i_17_n_0 ),
        .O(\instruction[1]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h6))
    \instruction[1]_i_26
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA888AAAAA))
    \instruction[1]_i_27
       (.I0(\instruction_reg[1]_i_48_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\instruction[23]_i_22_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hB88BBBBBBBBBBBBB))
    \instruction[1]_i_28
       (.I0(\instruction[1]_i_49_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\instruction[5]_i_6_n_0 ),
        .O(\instruction[1]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0044A28000011000))
    \instruction[1]_i_29
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFDFFFF7FFF7DFFF))
    \instruction[1]_i_3
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .O(\instruction[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000050010800018))
    \instruction[1]_i_30
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h8AAAAAAA8AAA8A8A))
    \instruction[1]_i_31
       (.I0(\instruction_reg[1]_i_50_n_0 ),
        .I1(\instruction[7]_i_17_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hBEFEFFBEFFBEEE5E))
    \instruction[1]_i_32
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[1]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hDB49A5FFEDFEFF7F))
    \instruction[1]_i_33
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[1]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF3FFFFFFBFEFF))
    \instruction[1]_i_34
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[1]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0800100000000800))
    \instruction[1]_i_35
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\instruction[23]_i_22_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[1]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0080008000100000))
    \instruction[1]_i_36
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[1]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h0000A40000000000))
    \instruction[1]_i_37
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[1]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hEFFFFFFFEFFF0000))
    \instruction[1]_i_38
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\instruction[1]_i_51_n_0 ),
        .O(\instruction[1]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hF5B5FFBFFFFBFBFF))
    \instruction[1]_i_39
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[1]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFD5EFDF0FFFFFD))
    \instruction[1]_i_40
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[1]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0000400038000008))
    \instruction[1]_i_41
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[1]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0000000018040400))
    \instruction[1]_i_42
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[1]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000004020004000))
    \instruction[1]_i_43
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[1]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFF9FF))
    \instruction[1]_i_44
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\instruction_reg[1]_i_52_n_0 ),
        .O(\instruction[1]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA2AAAAAAAAAA))
    \instruction[1]_i_45
       (.I0(\instruction_reg[1]_i_53_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[1]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFEF7FFFFFFF77FFE))
    \instruction[1]_i_46
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[1]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000002000102))
    \instruction[1]_i_47
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[1]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFF7FFFDFFDDDFFF))
    \instruction[1]_i_49
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[1]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFDBFFABFFFB5))
    \instruction[1]_i_51
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[1]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hF5FFF5FFF7FFE7BF))
    \instruction[1]_i_54
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[1]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEFEF7FFF7FEFF))
    \instruction[1]_i_55
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[1]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFC79FFFF37DE7))
    \instruction[1]_i_56
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[1]_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFE7FFF9E))
    \instruction[1]_i_57
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[1]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'h0004010109042290))
    \instruction[1]_i_58
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[1]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hD500D50080208000))
    \instruction[1]_i_59
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[1]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h7F907FDF3DFF7DFF))
    \instruction[1]_i_60
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[1]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFCBFF7))
    \instruction[1]_i_61
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[1]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDFFF7DDF7FDF))
    \instruction[1]_i_8
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFDFFDFFFEFF))
    \instruction[1]_i_9
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h808080FFFFFF80FF))
    \instruction[20]_i_1
       (.I0(\instruction[20]_i_2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\instruction[20]_i_3_n_0 ),
        .I3(\instruction[20]_i_4_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction[20]_i_5_n_0 ),
        .O(\instruction[20]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h02))
    \instruction[20]_i_10
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[20]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h3747347774477747))
    \instruction[20]_i_11
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[20]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000026))
    \instruction[20]_i_13
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\instruction[20]_i_20_n_0 ),
        .O(\instruction[20]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000036000000000))
    \instruction[20]_i_14
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\instruction[20]_i_21_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[20]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF7070000F707F707))
    \instruction[20]_i_15
       (.I0(\instruction[20]_i_22_n_0 ),
        .I1(\instruction[24]_i_15_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\instruction_reg[20]_i_23_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\instruction[20]_i_24_n_0 ),
        .O(\instruction[20]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h2EEE00002EEE2EEE))
    \instruction[20]_i_16
       (.I0(\instruction_reg[20]_i_25_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\instruction[20]_i_26_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\instruction[20]_i_27_n_0 ),
        .O(\instruction[20]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h37BFFFFC))
    \instruction[20]_i_17
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[20]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h048282A688000214))
    \instruction[20]_i_18
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[20]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h081B000C4206000C))
    \instruction[20]_i_19
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[20]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00D1FFFF00D10000))
    \instruction[20]_i_2
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\instruction[20]_i_6_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\instruction[20]_i_7_n_0 ),
        .O(\instruction[20]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[20]_i_20
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[20]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h7F))
    \instruction[20]_i_21
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[20]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h24))
    \instruction[20]_i_22
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[20]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h8000))
    \instruction[20]_i_24
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[20]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h000800D5F292F207))
    \instruction[20]_i_26
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[20]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h4000))
    \instruction[20]_i_27
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[20]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFE67FAAFFFA7))
    \instruction[20]_i_28
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[20]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hEFFFAFBFFFEBFEFF))
    \instruction[20]_i_29
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[20]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'hB))
    \instruction[20]_i_3
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h55DFFFDFFFDFFFDF))
    \instruction[20]_i_30
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[20]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h577F777FFF3FFF7F))
    \instruction[20]_i_31
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[20]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hA202A2A2A2A2A2A2))
    \instruction[20]_i_4
       (.I0(\instruction_reg[20]_i_8_n_0 ),
        .I1(\instruction[20]_i_9_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\instruction[25]_i_7_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\instruction[20]_i_10_n_0 ),
        .O(\instruction[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000008BFFFF))
    \instruction[20]_i_5
       (.I0(\instruction[20]_i_11_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\instruction_reg[20]_i_12_n_0 ),
        .I3(\instruction[20]_i_13_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\instruction[20]_i_14_n_0 ),
        .O(\instruction[20]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hEFEFFFFB))
    \instruction[20]_i_6
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC0100C0000000000))
    \instruction[20]_i_7
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[20]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00004041))
    \instruction[20]_i_9
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\instruction[20]_i_17_n_0 ),
        .O(\instruction[20]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5757F757F7F7F7F7))
    \instruction[21]_i_1
       (.I0(\instruction[21]_i_2_n_0 ),
        .I1(\instruction[21]_i_3_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[0] ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\instruction_reg[21]_i_4_n_0 ),
        .I5(\instruction_reg[21]_i_5_n_0 ),
        .O(\instruction[21]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000))
    \instruction[21]_i_12
       (.I0(\instruction[21]_i_29_n_0 ),
        .I1(\instruction[21]_i_30_n_0 ),
        .I2(\instruction[21]_i_31_n_0 ),
        .I3(\instruction[21]_i_32_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\instruction_reg[21]_i_33_n_0 ),
        .O(\instruction[21]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFBF3FBFFDBF3FBFF))
    \instruction[21]_i_14
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[21]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFAFFEFBFE))
    \instruction[21]_i_15
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[21]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00002E22))
    \instruction[21]_i_16
       (.I0(\instruction_reg[21]_i_36_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\instruction[21]_i_37_n_0 ),
        .I3(\instruction[21]_i_38_n_0 ),
        .I4(\instruction_reg[21]_i_39_n_0 ),
        .O(\instruction[21]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2222222))
    \instruction[21]_i_17
       (.I0(\instruction_reg[21]_i_40_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\instruction[21]_i_41_n_0 ),
        .I3(\instruction[21]_i_42_n_0 ),
        .I4(\instruction[21]_i_43_n_0 ),
        .I5(\instruction_reg[21]_i_44_n_0 ),
        .O(\instruction[21]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0212420400100000))
    \instruction[21]_i_18
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1205000812001000))
    \instruction[21]_i_19
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[21]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA8AAAAAA))
    \instruction[21]_i_2
       (.I0(\instruction[21]_i_6_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[2] ),
        .I3(\instruction[21]_i_7_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\instruction[21]_i_8_n_0 ),
        .O(\instruction[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000040FFFFFFFF))
    \instruction[21]_i_20
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep_n_0_[2] ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\instruction[21]_i_45_n_0 ),
        .I5(\instruction[21]_i_46_n_0 ),
        .O(\instruction[21]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8000BB0800000044))
    \instruction[21]_i_21
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[21]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000010100F0000))
    \instruction[21]_i_22
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[21]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCC0CCCCCCC4C4))
    \instruction[21]_i_23
       (.I0(\instruction[25]_i_11_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[21]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFBF5D6FDF67BBC))
    \instruction[21]_i_24
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[21]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hC66FDBBFDBF7EFFF))
    \instruction[21]_i_25
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[21]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hDBBFDF7FD76BBFF7))
    \instruction[21]_i_26
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h2168600604800120))
    \instruction[21]_i_27
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[21]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hE829944228004029))
    \instruction[21]_i_28
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[21]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h6))
    \instruction[21]_i_29
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[21]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004F40404))
    \instruction[21]_i_3
       (.I0(\instruction[21]_i_9_n_0 ),
        .I1(\instruction_reg[21]_i_10_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\instruction_reg[21]_i_11_n_0 ),
        .I4(\instruction[21]_i_12_n_0 ),
        .I5(\instruction_reg[21]_i_13_n_0 ),
        .O(\instruction[21]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[21]_i_30
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[21]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h0206))
    \instruction[21]_i_31
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFCF4FFF00FFFF4F))
    \instruction[21]_i_32
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[21]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0311A2104711A200))
    \instruction[21]_i_37
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[21]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEFFFFBBFEFFFE))
    \instruction[21]_i_38
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[21]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FFD0FFDD))
    \instruction[21]_i_41
       (.I0(\instruction[21]_i_59_n_0 ),
        .I1(\instruction[16]_i_11_n_0 ),
        .I2(\instruction[21]_i_60_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .I5(\instruction[21]_i_61_n_0 ),
        .O(\instruction[21]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h7F7FFFFFFFFF7FFF))
    \instruction[21]_i_42
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[21]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFDFF5DF))
    \instruction[21]_i_43
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_43_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[21]_i_45
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[21]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFDFFFFFF))
    \instruction[21]_i_46
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFEFDFFFEFB7FEBF7))
    \instruction[21]_i_47
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[21]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFF6BFFFFEBF7))
    \instruction[21]_i_48
       (.I0(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[21]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h8800880020002001))
    \instruction[21]_i_49
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[21]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0088008004560000))
    \instruction[21]_i_50
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[21]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000020))
    \instruction[21]_i_51
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[21]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00AA000055554200))
    \instruction[21]_i_52
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[21]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hEFDFF66DFEEFDFFF))
    \instruction[21]_i_53
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[21]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDFDEF7FF6D6FD))
    \instruction[21]_i_54
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[21]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hA410200040841060))
    \instruction[21]_i_55
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[21]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h4914400040008440))
    \instruction[21]_i_56
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDEDFFFF7EFED7))
    \instruction[21]_i_57
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[21]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hEFFEFEFBEFEFFFBF))
    \instruction[21]_i_58
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[21]_i_58_n_0 ));
  LUT3 #(
    .INIT(8'h9A))
    \instruction[21]_i_59
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h55555555F5F7FDFF))
    \instruction[21]_i_6
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\instruction[21]_i_18_n_0 ),
        .I4(\instruction[21]_i_19_n_0 ),
        .I5(\instruction[21]_i_20_n_0 ),
        .O(\instruction[21]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[21]_i_60
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .O(\instruction[21]_i_60_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[21]_i_61
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h3029900094402004))
    \instruction[21]_i_62
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[21]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h5442299421804001))
    \instruction[21]_i_63
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[21]_i_63_n_0 ));
  LUT2 #(
    .INIT(4'h8))
    \instruction[21]_i_7
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[21]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[21]_i_8
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[21]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222F0002222F0FF))
    \instruction[21]_i_9
       (.I0(\instruction[21]_i_21_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\instruction[21]_i_22_n_0 ),
        .I3(\instruction[21]_i_23_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\instruction[21]_i_24_n_0 ),
        .O(\instruction[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00008000FFFFFFFF))
    \instruction[22]_i_1
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[9] ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction[22]_i_2_n_0 ),
        .O(\instruction[22]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFBFFFBFFBBDDEF))
    \instruction[22]_i_10
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\program_counter_reg_rep_n_0_[1] ),
        .O(\instruction[22]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h80AF40004050C000))
    \instruction[22]_i_11
       (.I0(\program_counter_reg_rep_n_0_[0] ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[9] ),
        .I5(\program_counter_reg_rep_n_0_[1] ),
        .O(\instruction[22]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF))
    \instruction[22]_i_12
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep_n_0_[1] ),
        .O(\instruction[22]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h06000000))
    \instruction[22]_i_13
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep_n_0_[0] ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[9] ),
        .O(\instruction[22]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h1FFFFFFF1FFF0000))
    \instruction[22]_i_2
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep_n_0_[9] ),
        .I3(\instruction[22]_i_3_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\instruction[22]_i_4_n_0 ),
        .O(\instruction[22]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h01000000FFFFFFFF))
    \instruction[22]_i_3
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep_n_0_[0] ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\instruction_reg[22]_i_5_n_0 ),
        .O(\instruction[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFF7FF0000))
    \instruction[22]_i_4
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\instruction[22]_i_6_n_0 ),
        .I3(\instruction[22]_i_7_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\instruction[22]_i_8_n_0 ),
        .O(\instruction[22]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[22]_i_6
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[22]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEA404044406240EA))
    \instruction[22]_i_7
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[0] ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\program_counter_reg_rep_n_0_[9] ),
        .O(\instruction[22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4444FFFC7774FFFC))
    \instruction[22]_i_8
       (.I0(\instruction[22]_i_11_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[9] ),
        .I3(\instruction[22]_i_12_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\instruction[22]_i_13_n_0 ),
        .O(\instruction[22]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBD4DFFFF))
    \instruction[22]_i_9
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep_n_0_[0] ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[22]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFDF55DFFFDFFFDF))
    \instruction[23]_i_1
       (.I0(\instruction_reg[23]_i_2_n_0 ),
        .I1(\instruction[23]_i_3_n_0 ),
        .I2(\instruction_reg[23]_i_4_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction_reg[23]_i_5_n_0 ),
        .I5(\instruction_reg[23]_i_6_n_0 ),
        .O(\instruction[23]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF5FFFFF5F77F7F7F))
    \instruction[23]_i_11
       (.I0(\instruction[23]_i_22_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[23]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h888888B8B8B888B8))
    \instruction[23]_i_12
       (.I0(\instruction[23]_i_23_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[23]_i_24_n_0 ),
        .I3(\instruction[23]_i_25_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\instruction[23]_i_26_n_0 ),
        .O(\instruction[23]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h8000808080808080))
    \instruction[23]_i_13
       (.I0(\instruction_reg[23]_i_27_n_0 ),
        .I1(\instruction[23]_i_28_n_0 ),
        .I2(\instruction[23]_i_29_n_0 ),
        .I3(\instruction[23]_i_30_n_0 ),
        .I4(\instruction[23]_i_31_n_0 ),
        .I5(\instruction[23]_i_32_n_0 ),
        .O(\instruction[23]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8BB88))
    \instruction[23]_i_14
       (.I0(\instruction_reg[23]_i_33_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[23]_i_34_n_0 ),
        .I3(\instruction[23]_i_35_n_0 ),
        .I4(\instruction[23]_i_36_n_0 ),
        .O(\instruction[23]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAC00ACFFACFFACFF))
    \instruction[23]_i_15
       (.I0(\instruction[23]_i_37_n_0 ),
        .I1(\instruction[23]_i_38_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\instruction[23]_i_39_n_0 ),
        .I5(\instruction_reg[23]_i_40_n_0 ),
        .O(\instruction[23]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF))
    \instruction[23]_i_16
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[23]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBB8BBBBBBBBBB))
    \instruction[23]_i_17
       (.I0(\instruction[23]_i_41_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\instruction[25]_i_9_n_0 ),
        .O(\instruction[23]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0002020002000000))
    \instruction[23]_i_18
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[23]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0080FFFF00800000))
    \instruction[23]_i_19
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\instruction[23]_i_42_n_0 ),
        .O(\instruction[23]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFF7F7F7FBFFFBFF))
    \instruction[23]_i_20
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[23]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h777FFFDFFF0FFFFF))
    \instruction[23]_i_21
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[23]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[23]_i_22
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[23]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA2AAA2AAAAAA))
    \instruction[23]_i_23
       (.I0(\instruction_reg[23]_i_43_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hDBBDDFFBFFFFBDF7))
    \instruction[23]_i_24
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0040099009940020))
    \instruction[23]_i_25
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[23]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000A58181))
    \instruction[23]_i_26
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[23]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h5FFFFFFFFFDFFF7D))
    \instruction[23]_i_28
       (.I0(\instruction[23]_i_46_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[23]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF))
    \instruction[23]_i_29
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\instruction[23]_i_47_n_0 ),
        .O(\instruction[23]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h101010FFFFFF10FF))
    \instruction[23]_i_3
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\instruction[23]_i_9_n_0 ),
        .I3(\instruction_reg[23]_i_10_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\instruction[23]_i_11_n_0 ),
        .O(\instruction[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[23]_i_30
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[23]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h40))
    \instruction[23]_i_31
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[23]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[23]_i_32
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[23]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h1100110010FF1000))
    \instruction[23]_i_34
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[23]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h249212494B24A492))
    \instruction[23]_i_35
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[23]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h2022AAAA))
    \instruction[23]_i_36
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[23]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000E2E200))
    \instruction[23]_i_37
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[23]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hE118826118866118))
    \instruction[23]_i_38
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[23]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hDBBDD77FFFFFBFF6))
    \instruction[23]_i_39
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h57FFFFFFFFFFFFEF))
    \instruction[23]_i_41
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[23]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h8380000C80800000))
    \instruction[23]_i_42
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[23]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[23]_i_46
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[23]_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[23]_i_47
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[23]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0502021010052502))
    \instruction[23]_i_48
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[23]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hAABA449201014924))
    \instruction[23]_i_49
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFEDB2FB6FB7))
    \instruction[23]_i_50
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000FBFE7FDFFFEF))
    \instruction[23]_i_51
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hEFFDFDDADAEFEFFD))
    \instruction[23]_i_52
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[23]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hFDFEFEF7F7FDB9BE))
    \instruction[23]_i_53
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFEEDDBB6DBF66DDB))
    \instruction[23]_i_54
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFD8EDEE7E7797DDF))
    \instruction[23]_i_55
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[23]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFBFF0BFF0BFFF))
    \instruction[23]_i_56
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[23]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF0035FFBCFF))
    \instruction[23]_i_57
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[23]_i_57_n_0 ));
  LUT5 #(
    .INIT(32'hFFF75DFF))
    \instruction[23]_i_7
       (.I0(\instruction[23]_i_18_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[23]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h2FBEFFFF))
    \instruction[23]_i_8
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\instruction[23]_i_19_n_0 ),
        .O(\instruction[23]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h0080))
    \instruction[23]_i_9
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[23]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF777FFFF))
    \instruction[24]_i_1
       (.I0(\instruction[24]_i_2_n_0 ),
        .I1(\instruction_reg[24]_i_3_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\instruction_reg[24]_i_4_n_0 ),
        .I4(\instruction_reg[24]_i_5_n_0 ),
        .O(\instruction[24]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h20FF2902))
    \instruction[24]_i_10
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[24]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h2E22000000000000))
    \instruction[24]_i_11
       (.I0(\instruction[24]_i_18_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\instruction_reg[24]_i_19_n_0 ),
        .I3(\instruction_reg[24]_i_20_n_0 ),
        .I4(\instruction[24]_i_21_n_0 ),
        .I5(\instruction[24]_i_22_n_0 ),
        .O(\instruction[24]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00E2E2E200000000))
    \instruction[24]_i_12
       (.I0(\instruction[24]_i_23_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\instruction[24]_i_24_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\instruction_reg[24]_i_25_n_0 ),
        .I5(\instruction[24]_i_26_n_0 ),
        .O(\instruction[24]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4FFF4AAAAAAAA))
    \instruction[24]_i_13
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\instruction[24]_i_27_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[24]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAA8082AAAA80A280))
    \instruction[24]_i_14
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[24]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0040))
    \instruction[24]_i_15
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[24]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hD775555555555555))
    \instruction[24]_i_16
       (.I0(\instruction[24]_i_28_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\instruction[24]_i_29_n_0 ),
        .I5(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[24]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100))
    \instruction[24]_i_17
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\instruction[24]_i_30_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .O(\instruction[24]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040737F7F))
    \instruction[24]_i_18
       (.I0(\instruction[24]_i_31_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\instruction[24]_i_32_n_0 ),
        .I5(\instruction[24]_i_33_n_0 ),
        .O(\instruction[24]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF7FFFFF7F7FF))
    \instruction[24]_i_2
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\instruction[24]_i_6_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFE0EFEFEFEFEFEFE))
    \instruction[24]_i_21
       (.I0(\instruction[24]_i_38_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[24]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h3FFF3FFF0F7FBF7F))
    \instruction[24]_i_22
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[24]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h000000E2E2E200E2))
    \instruction[24]_i_23
       (.I0(\instruction[24]_i_39_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\instruction[24]_i_40_n_0 ),
        .I3(\instruction_reg[24]_i_41_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\instruction[24]_i_42_n_0 ),
        .O(\instruction[24]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h000000E2E2E200E2))
    \instruction[24]_i_24
       (.I0(\instruction[24]_i_43_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[24]_i_44_n_0 ),
        .I3(\instruction_reg[24]_i_45_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\instruction[24]_i_46_n_0 ),
        .O(\instruction[24]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF6FFFFFF))
    \instruction[24]_i_26
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .O(\instruction[24]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[24]_i_27
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[24]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFFFABFF))
    \instruction[24]_i_28
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\instruction[19]_i_18_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\instruction[24]_i_49_n_0 ),
        .O(\instruction[24]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[24]_i_29
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[24]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[24]_i_30
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[24]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'h0000C088))
    \instruction[24]_i_31
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[24]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h034CC04C004CC04C))
    \instruction[24]_i_32
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[24]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888))
    \instruction[24]_i_33
       (.I0(\instruction[24]_i_50_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\instruction[24]_i_51_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\instruction[24]_i_52_n_0 ),
        .O(\instruction[24]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h9000009000000010))
    \instruction[24]_i_34
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\instruction[25]_i_8_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[24]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFB400000000))
    \instruction[24]_i_35
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .O(\instruction[24]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h77BDBF6F6BD7DFBF))
    \instruction[24]_i_36
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[24]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h6F6B6FDFD6BFBF6F))
    \instruction[24]_i_37
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[24]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFF33CFFFFF77FFF))
    \instruction[24]_i_38
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[24]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hBFB797FB77FBFBFF))
    \instruction[24]_i_39
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .O(\instruction[24]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hCDEB6BDEDEFFBDFF))
    \instruction[24]_i_40
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[24]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h4004400440044007))
    \instruction[24]_i_42
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[24]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h4D6B6FDFD6BFBFEF))
    \instruction[24]_i_43
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[24]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hBBBDD77FD66BBFFF))
    \instruction[24]_i_44
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[24]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h28280000282800FC))
    \instruction[24]_i_46
       (.I0(\instruction[24]_i_57_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[24]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'h00000880))
    \instruction[24]_i_47
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[24]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h30C030AF000000AA))
    \instruction[24]_i_48
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[24]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA00003A0A))
    \instruction[24]_i_49
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[24]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h4D24499249922449))
    \instruction[24]_i_50
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[24]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0050005018218080))
    \instruction[24]_i_51
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[24]_i_51_n_0 ));
  LUT5 #(
    .INIT(32'h82080820))
    \instruction[24]_i_52
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[24]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002400))
    \instruction[24]_i_53
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[24]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h4100000000824100))
    \instruction[24]_i_54
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[24]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000041800080000))
    \instruction[24]_i_55
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .O(\instruction[24]_i_55_n_0 ));
  LUT5 #(
    .INIT(32'h04000000))
    \instruction[24]_i_56
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[24]_i_56_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[24]_i_57
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[24]_i_57_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[24]_i_6
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[24]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h7777077777777777))
    \instruction[24]_i_7
       (.I0(\instruction[24]_i_13_n_0 ),
        .I1(\instruction[24]_i_14_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\instruction[24]_i_15_n_0 ),
        .O(\instruction[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4747474747470047))
    \instruction[24]_i_8
       (.I0(\instruction[24]_i_16_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\instruction[24]_i_17_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\instruction[21]_i_8_n_0 ),
        .I5(\instruction[24]_i_6_n_0 ),
        .O(\instruction[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h3170315000080042))
    \instruction[24]_i_9
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[24]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFDF55DFFFDFFFDF))
    \instruction[25]_i_1
       (.I0(\instruction[25]_i_2_n_0 ),
        .I1(\instruction[25]_i_3_n_0 ),
        .I2(\instruction_reg[25]_i_4_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction[25]_i_5_n_0 ),
        .I5(\instruction[25]_i_6_n_0 ),
        .O(\instruction[25]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8))
    \instruction[25]_i_10
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[25]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[25]_i_11
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[25]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAA2AAAAA))
    \instruction[25]_i_12
       (.I0(\instruction_reg[25]_i_20_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[25]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000000000407F4F7))
    \instruction[25]_i_13
       (.I0(\instruction[25]_i_21_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\instruction[25]_i_22_n_0 ),
        .I3(\instruction[25]_i_23_n_0 ),
        .I4(\instruction[25]_i_24_n_0 ),
        .I5(\instruction[25]_i_25_n_0 ),
        .O(\instruction[25]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[25]_i_14
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[25]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[25]_i_15
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[25]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA8AAAAAAA))
    \instruction[25]_i_16
       (.I0(\instruction_reg[25]_i_26_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[25]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hEEEAEEEE222A2222))
    \instruction[25]_i_17
       (.I0(\instruction[25]_i_27_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\instruction[25]_i_28_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\instruction[25]_i_29_n_0 ),
        .O(\instruction[25]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF))
    \instruction[25]_i_18
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[25]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFFFFFFFF))
    \instruction[25]_i_2
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\instruction[25]_i_7_n_0 ),
        .I2(\instruction[25]_i_8_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\instruction[25]_i_9_n_0 ),
        .O(\instruction[25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0881166816688116))
    \instruction[25]_i_21
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[25]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAA800000000))
    \instruction[25]_i_22
       (.I0(\instruction[25]_i_35_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\instruction[25]_i_28_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[25]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h6449499292242448))
    \instruction[25]_i_23
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[2] ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[25]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0014080000000222))
    \instruction[25]_i_24
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[25]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000))
    \instruction[25]_i_25
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[4]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[25]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hEBD6DEBDD6BDBD6B))
    \instruction[25]_i_27
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[25]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'hB))
    \instruction[25]_i_28
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[25]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFBFFB))
    \instruction[25]_i_29
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[25]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hC000000000001000))
    \instruction[25]_i_3
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\instruction[25]_i_10_n_0 ),
        .I3(\instruction[25]_i_11_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h7777F7FF5555F5F5))
    \instruction[25]_i_30
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\instruction[25]_i_38_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\instruction[25]_i_39_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[25]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEFEBFFFFFFEBF))
    \instruction[25]_i_35
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[25]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hBF76FEE9EBBFBFF4))
    \instruction[25]_i_36
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[25]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBFFD6EB46E6ED))
    \instruction[25]_i_37
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[25]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hFD))
    \instruction[25]_i_38
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .O(\instruction[25]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'hB))
    \instruction[25]_i_39
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .O(\instruction[25]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h00002804))
    \instruction[25]_i_40
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[25]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'h40040004))
    \instruction[25]_i_41
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[25]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0229904294422994))
    \instruction[25]_i_42
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[25]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h044229942D944229))
    \instruction[25]_i_43
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[25]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hBBB66DDB6DDBB66D))
    \instruction[25]_i_44
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[25]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hB66DDBB6DBF66DDB))
    \instruction[25]_i_45
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[4]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[25]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFE5FFF5EBAFEFFFE))
    \instruction[25]_i_46
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[25]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFBABFFFFEFFEFFFB))
    \instruction[25]_i_47
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[4]_rep_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[25]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00E0000000000020))
    \instruction[25]_i_5
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\instruction[25]_i_14_n_0 ),
        .I3(\instruction[25]_i_15_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[25]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB800B800B8FFB800))
    \instruction[25]_i_6
       (.I0(\instruction[25]_i_16_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\instruction[25]_i_17_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\instruction[25]_i_18_n_0 ),
        .I5(\instruction_reg[25]_i_19_n_0 ),
        .O(\instruction[25]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[25]_i_7
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[25]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[25]_i_8
       (.I0(\program_counter_reg_rep[4]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[25]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[25]_i_9
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[25]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D1DFFFFFF1DFF))
    \instruction[26]_i_1
       (.I0(\instruction[26]_i_2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\instruction[26]_i_3_n_0 ),
        .I3(\instruction[26]_i_4_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction[26]_i_5_n_0 ),
        .O(\instruction[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000))
    \instruction[26]_i_11
       (.I0(\instruction[26]_i_17_n_0 ),
        .I1(\instruction[25]_i_9_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[26]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0FFFFFFFEFFFF))
    \instruction[26]_i_12
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\instruction[25]_i_7_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\instruction[26]_i_18_n_0 ),
        .O(\instruction[26]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h07000FFF07FF0FFF))
    \instruction[26]_i_13
       (.I0(\instruction[26]_i_19_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[26]_i_20_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\instruction_reg[26]_i_21_n_0 ),
        .O(\instruction[26]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8121000080204040))
    \instruction[26]_i_14
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[26]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hC422008881002301))
    \instruction[26]_i_15
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep_n_0_[3] ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[26]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h080A140249995444))
    \instruction[26]_i_16
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[3] ),
        .O(\instruction[26]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[26]_i_17
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[26]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h8000))
    \instruction[26]_i_18
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[26]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100602))
    \instruction[26]_i_19
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[5]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[26]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h57F7F7F7))
    \instruction[26]_i_2
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\instruction[26]_i_6_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8888F8F8FF88F8F8))
    \instruction[26]_i_20
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\instruction[26]_i_18_n_0 ),
        .I2(\instruction[26]_i_22_n_0 ),
        .I3(\instruction[26]_i_23_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[26]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000240000000000))
    \instruction[26]_i_22
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\instruction[25]_i_9_n_0 ),
        .O(\instruction[26]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0C380C000C000C00))
    \instruction[26]_i_23
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[26]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h00000188))
    \instruction[26]_i_24
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[26]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h8AA080808A8080A2))
    \instruction[26]_i_25
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[26]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hF757F7F7F7F7F7F7))
    \instruction[26]_i_3
       (.I0(\instruction[26]_i_7_n_0 ),
        .I1(\instruction[26]_i_8_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep_n_0 ),
        .O(\instruction[26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h470047FF00000000))
    \instruction[26]_i_4
       (.I0(\instruction[26]_i_9_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\instruction_reg[26]_i_10_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\instruction[26]_i_11_n_0 ),
        .I5(\instruction[26]_i_12_n_0 ),
        .O(\instruction[26]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h2AA8A2A2AAAAAAAA))
    \instruction[26]_i_5
       (.I0(\instruction[26]_i_13_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep_n_0_[7] ),
        .I4(\program_counter_reg_rep[5]_rep_n_0 ),
        .I5(\instruction[26]_i_14_n_0 ),
        .O(\instruction[26]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00000040))
    \instruction[26]_i_6
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[26]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hA202))
    \instruction[26]_i_7
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[5]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[26]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hD0D0C000000F0000))
    \instruction[26]_i_8
       (.I0(\program_counter_reg_rep[5]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h020C020C07000207))
    \instruction[26]_i_9
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[5]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[26]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000080FFFFFFFF))
    \instruction[27]_i_1
       (.I0(\program_counter_reg_rep_n_0_[0] ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\instruction[27]_i_2_n_0 ),
        .I5(\instruction_reg[27]_i_3_n_0 ),
        .O(\instruction[27]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0282FFFF02820000))
    \instruction[27]_i_10
       (.I0(\program_counter_reg_rep_n_0_[0] ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\instruction[27]_i_13_n_0 ),
        .O(\instruction[27]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4400440040104900))
    \instruction[27]_i_11
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[6]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[27]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h200022004D312200))
    \instruction[27]_i_13
       (.I0(\program_counter_reg_rep_n_0_[0] ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[27]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBFBFFFFFFFBFF))
    \instruction[27]_i_14
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep_n_0_[7] ),
        .O(\instruction[27]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h7F7F7FFFFFFFF6FF))
    \instruction[27]_i_15
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[7] ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[27]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[27]_i_2
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7))
    \instruction[27]_i_4
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\instruction[27]_i_6_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[0] ),
        .I3(\instruction[27]_i_7_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\instruction[27]_i_8_n_0 ),
        .O(\instruction[27]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h2AAAAAAA))
    \instruction[27]_i_5
       (.I0(\instruction[27]_i_9_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0033004000000340))
    \instruction[27]_i_6
       (.I0(\program_counter_reg_rep[6]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep_n_0_[7] ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000070000004))
    \instruction[27]_i_7
       (.I0(\program_counter_reg_rep_n_0_[7] ),
        .I1(\program_counter_reg_rep[6]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h001080B0808F8080))
    \instruction[27]_i_8
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\instruction[25]_i_28_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\program_counter_reg_rep_n_0_[1] ),
        .O(\instruction[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4F7F7F7F4F7F4C4C))
    \instruction[27]_i_9
       (.I0(\instruction[27]_i_10_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\instruction[27]_i_11_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction_reg[27]_i_12_n_0 ),
        .O(\instruction[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFDF55DFFFDFFFDF))
    \instruction[2]_i_1
       (.I0(\instruction_reg[2]_i_2_n_0 ),
        .I1(\instruction[2]_i_3_n_0 ),
        .I2(\instruction_reg[2]_i_4_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction_reg[2]_i_5_n_0 ),
        .I5(\instruction[2]_i_6_n_0 ),
        .O(\instruction[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000800))
    \instruction[2]_i_10
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFF7FFF))
    \instruction[2]_i_11
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\instruction[2]_i_26_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00E2E2E2E2E2E2E2))
    \instruction[2]_i_12
       (.I0(\instruction[2]_i_27_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction_reg[2]_i_28_n_0 ),
        .I3(\instruction[2]_i_29_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\instruction[7]_i_11_n_0 ),
        .O(\instruction[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h0000440C))
    \instruction[2]_i_13
       (.I0(\instruction_reg[2]_i_30_n_0 ),
        .I1(\instruction_reg[2]_i_31_n_0 ),
        .I2(\instruction[2]_i_32_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\instruction[2]_i_33_n_0 ),
        .O(\instruction[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000004000200000))
    \instruction[2]_i_14
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\instruction[3]_i_23_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0808100200000000))
    \instruction[2]_i_15
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\instruction[6]_i_13_n_0 ),
        .O(\instruction[2]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hF7))
    \instruction[2]_i_17
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[2]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[2]_i_18
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000018000220))
    \instruction[2]_i_20
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[2]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00881480A0000000))
    \instruction[2]_i_21
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[2]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h02))
    \instruction[2]_i_22
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[2]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h80))
    \instruction[2]_i_23
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[2]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hBBFFEEFFFFFEFFFF))
    \instruction[2]_i_24
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[2]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h04000000))
    \instruction[2]_i_25
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[2]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[2]_i_26
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[2]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAABA0000AA8A))
    \instruction[2]_i_27
       (.I0(\instruction[2]_i_39_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I5(\instruction[2]_i_40_n_0 ),
        .O(\instruction[2]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[2]_i_29
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[2]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0FFF4FF))
    \instruction[2]_i_3
       (.I0(\instruction[2]_i_9_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\instruction[2]_i_10_n_0 ),
        .I3(\instruction[2]_i_11_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h08FF080008000800))
    \instruction[2]_i_32
       (.I0(\instruction[17]_i_25_n_0 ),
        .I1(\instruction[23]_i_22_n_0 ),
        .I2(\instruction[4]_i_29_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\instruction[7]_i_11_n_0 ),
        .O(\instruction[2]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0024410000000000))
    \instruction[2]_i_33
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\instruction[2]_i_47_n_0 ),
        .O(\instruction[2]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hA8AA8A88AAAAAAAA))
    \instruction[2]_i_34
       (.I0(\instruction_reg[2]_i_48_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\instruction[2]_i_49_n_0 ),
        .O(\instruction[2]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hF5FF77E7FFFFFFFF))
    \instruction[2]_i_35
       (.I0(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\instruction[2]_i_50_n_0 ),
        .O(\instruction[2]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hD5555555))
    \instruction[2]_i_36
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[2]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFEBF93D00DEFB4B))
    \instruction[2]_i_39
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[2]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFBBEFB7FF6DEBFB))
    \instruction[2]_i_40
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[2]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFEFFEFF))
    \instruction[2]_i_41
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[2]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hDFF01FFFDFFF1FFF))
    \instruction[2]_i_42
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[2]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h043402011C1C0598))
    \instruction[2]_i_43
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[2]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h4008170820282128))
    \instruction[2]_i_44
       (.I0(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[2]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hBFBFBFFFFFFFBFFF))
    \instruction[2]_i_45
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[2]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFF7FFFFDFFE7))
    \instruction[2]_i_46
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[2]_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[2]_i_47
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[2]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h24))
    \instruction[2]_i_49
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[2]_i_49_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[2]_i_50
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[2]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hF6FFFFF6DFDFFFFE))
    \instruction[2]_i_51
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[2]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hBBFFBFFFB3FFBFB3))
    \instruction[2]_i_52
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[2]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hFFAFFEEFEFFBFFFF))
    \instruction[2]_i_53
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[2]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h9F9E9F97009FFFF3))
    \instruction[2]_i_54
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[2]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFFF8FFFFAFAEDF3D))
    \instruction[2]_i_55
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[2]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFEF85FFEFFFFBBB7))
    \instruction[2]_i_56
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[2]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hAA8AFFFFAA8A0000))
    \instruction[2]_i_6
       (.I0(\instruction_reg[2]_i_16_n_0 ),
        .I1(\instruction[2]_i_17_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\instruction[2]_i_18_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\instruction_reg[2]_i_19_n_0 ),
        .O(\instruction[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4F7F40704F7F4F7F))
    \instruction[2]_i_7
       (.I0(\instruction[2]_i_20_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\instruction[2]_i_21_n_0 ),
        .I4(\instruction[7]_i_17_n_0 ),
        .I5(\instruction[18]_i_34_n_0 ),
        .O(\instruction[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7F7070707F707F7F))
    \instruction[2]_i_8
       (.I0(\instruction[2]_i_22_n_0 ),
        .I1(\instruction[2]_i_23_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\instruction[2]_i_24_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I5(\instruction[2]_i_25_n_0 ),
        .O(\instruction[2]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFB7FFD))
    \instruction[2]_i_9
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .O(\instruction[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBFBFFFFFFFBFF))
    \instruction[3]_i_1
       (.I0(\instruction[3]_i_2_n_0 ),
        .I1(\instruction_reg[3]_i_3_n_0 ),
        .I2(\instruction[3]_i_4_n_0 ),
        .I3(\instruction_reg[3]_i_5_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction[3]_i_6_n_0 ),
        .O(\instruction[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8))
    \instruction[3]_i_10
       (.I0(\instruction_reg[3]_i_24_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\instruction[2]_i_18_n_0 ),
        .O(\instruction[3]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100))
    \instruction[3]_i_11
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF6EFFFFFFFFFF))
    \instruction[3]_i_12
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\instruction[26]_i_17_n_0 ),
        .O(\instruction[3]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000000001105FFFF))
    \instruction[3]_i_15
       (.I0(\instruction[3]_i_29_n_0 ),
        .I1(\instruction[3]_i_30_n_0 ),
        .I2(\instruction[3]_i_31_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\instruction[3]_i_32_n_0 ),
        .O(\instruction[3]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000000E2E2E200E2))
    \instruction[3]_i_16
       (.I0(\instruction[3]_i_33_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\instruction[3]_i_34_n_0 ),
        .I3(\instruction[3]_i_35_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\instruction[3]_i_36_n_0 ),
        .O(\instruction[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFBFFEFFBFBFF))
    \instruction[3]_i_19
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hB88888B8888888B8))
    \instruction[3]_i_2
       (.I0(\instruction[3]_i_7_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\instruction[3]_i_8_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8083000000000000))
    \instruction[3]_i_20
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEFFFFFFFFFAFF))
    \instruction[3]_i_21
       (.I0(\instruction[3]_i_41_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \instruction[3]_i_23
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[3]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hEBFF5FFFFF7FFFF7))
    \instruction[3]_i_25
       (.I0(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[3]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFBFFBFFEFFFF))
    \instruction[3]_i_26
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000101010621500))
    \instruction[3]_i_27
       (.I0(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[3]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0000100410010088))
    \instruction[3]_i_28
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h08000000FFFFFFFF))
    \instruction[3]_i_29
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\instruction[3]_i_46_n_0 ),
        .O(\instruction[3]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h373C8844C4C80000))
    \instruction[3]_i_30
       (.I0(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h8091001120200100))
    \instruction[3]_i_31
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBFBBBBBFB))
    \instruction[3]_i_32
       (.I0(\instruction[3]_i_47_n_0 ),
        .I1(\instruction[3]_i_48_n_0 ),
        .I2(\instruction[3]_i_49_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h000000005F5FD5DF))
    \instruction[3]_i_33
       (.I0(\instruction[3]_i_50_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\instruction[3]_i_51_n_0 ),
        .O(\instruction[3]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAAAAAAAAAAAAA))
    \instruction[3]_i_34
       (.I0(\instruction_reg[3]_i_52_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0334884400008800))
    \instruction[3]_i_35
       (.I0(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[3]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000006101))
    \instruction[3]_i_36
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h0000F404))
    \instruction[3]_i_37
       (.I0(\instruction_reg[3]_i_53_n_0 ),
        .I1(\instruction[3]_i_54_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\instruction[3]_i_55_n_0 ),
        .I4(\instruction_reg[3]_i_56_n_0 ),
        .O(\instruction[3]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0000E200E200E200))
    \instruction[3]_i_38
       (.I0(\instruction_reg[3]_i_57_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\instruction[3]_i_58_n_0 ),
        .I3(\instruction_reg[3]_i_59_n_0 ),
        .I4(\instruction[3]_i_60_n_0 ),
        .I5(\instruction[3]_i_61_n_0 ),
        .O(\instruction[3]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF6EFFFFFFFF))
    \instruction[3]_i_39
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[3]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hBFBFFF3F))
    \instruction[3]_i_4
       (.I0(\instruction[3]_i_11_n_0 ),
        .I1(\instruction[3]_i_12_n_0 ),
        .I2(\instruction_reg[3]_i_13_n_0 ),
        .I3(\instruction_reg[3]_i_14_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8))
    \instruction[3]_i_40
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[3]_i_40_n_0 ));
  LUT2 #(
    .INIT(4'hB))
    \instruction[3]_i_41
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h2BFFB9D66FFFF5D7))
    \instruction[3]_i_42
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[3]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFF9FFFAFFFDFF9BF))
    \instruction[3]_i_43
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h007DFF7D00000000))
    \instruction[3]_i_44
       (.I0(\instruction[3]_i_62_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\instruction[3]_i_63_n_0 ),
        .I5(\instruction[3]_i_64_n_0 ),
        .O(\instruction[3]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAA2AAAAA))
    \instruction[3]_i_45
       (.I0(\instruction_reg[3]_i_65_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFDFEDDEEFFEF))
    \instruction[3]_i_46
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[3]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0044001100F40F11))
    \instruction[3]_i_47
       (.I0(\instruction[3]_i_66_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\instruction[3]_i_67_n_0 ),
        .O(\instruction[3]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFFFFFFFDFF5))
    \instruction[3]_i_48
       (.I0(\instruction[3]_i_68_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[3]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'h45406242))
    \instruction[3]_i_49
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[3]_i_49_n_0 ));
  LUT5 #(
    .INIT(32'h2244E24F))
    \instruction[3]_i_50
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[3]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h420000004A004202))
    \instruction[3]_i_51
       (.I0(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[3]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hABFFFFFFFFFFFFBF))
    \instruction[3]_i_54
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[3]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC000004440444))
    \instruction[3]_i_55
       (.I0(\instruction[3]_i_73_n_0 ),
        .I1(\instruction[3]_i_74_n_0 ),
        .I2(\instruction[3]_i_75_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\instruction[24]_i_6_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[3]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hEB5F5DEFFFF5F7FF))
    \instruction[3]_i_58
       (.I0(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[3]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h80808A8000000000))
    \instruction[3]_i_6
       (.I0(\instruction_reg[3]_i_17_n_0 ),
        .I1(\instruction_reg[3]_i_18_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\instruction[3]_i_19_n_0 ),
        .I4(\instruction[3]_i_20_n_0 ),
        .I5(\instruction[3]_i_21_n_0 ),
        .O(\instruction[3]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h04))
    \instruction[3]_i_60
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[3]_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h24))
    \instruction[3]_i_61
       (.I0(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[3]_i_61_n_0 ));
  LUT5 #(
    .INIT(32'h05056640))
    \instruction[3]_i_62
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[3]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000E00000))
    \instruction[3]_i_63
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[3]_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFFFFFDFFFFF3))
    \instruction[3]_i_64
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[3]_i_64_n_0 ));
  LUT3 #(
    .INIT(8'hEF))
    \instruction[3]_i_66
       (.I0(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[3]_i_66_n_0 ));
  LUT3 #(
    .INIT(8'hFE))
    \instruction[3]_i_67
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[3]_i_67_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[3]_i_68
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[3]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hC383FB8E3E30CFFF))
    \instruction[3]_i_69
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h0000000089040000))
    \instruction[3]_i_7
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFBFFFFFCFFFF0))
    \instruction[3]_i_70
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[6] ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0000822020349422))
    \instruction[3]_i_71
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .O(\instruction[3]_i_71_n_0 ));
  LUT5 #(
    .INIT(32'hA9208209))
    \instruction[3]_i_72
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[3]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h4300120041000055))
    \instruction[3]_i_73
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hB9F7FBB7FD5FF9BF))
    \instruction[3]_i_74
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[3]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'h04))
    \instruction[3]_i_75
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[3]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400200))
    \instruction[3]_i_76
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[3]_i_76_n_0 ));
  LUT5 #(
    .INIT(32'h00002410))
    \instruction[3]_i_77
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[3]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEF7F7))
    \instruction[3]_i_78
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[6] ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[3]_i_78_n_0 ));
  LUT6 #(
    .INIT(64'hEFFFFFFFFEFEEF5F))
    \instruction[3]_i_79
       (.I0(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[6] ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[3]_i_79_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004204020))
    \instruction[3]_i_8
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[6] ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFF7AEDFFFA7FFDD))
    \instruction[3]_i_80
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[6] ),
        .O(\instruction[3]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hB7BFFFD7BFFFFADF))
    \instruction[3]_i_81
       (.I0(\program_counter_reg_rep_n_0_[6] ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep_n_0 ),
        .O(\instruction[3]_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEFFFEFFFFFFFB))
    \instruction[3]_i_82
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDFFFDFFFFFFFD))
    \instruction[3]_i_83
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .O(\instruction[3]_i_83_n_0 ));
  LUT6 #(
    .INIT(64'hEAEEEEEEEEEEEEEE))
    \instruction[3]_i_9
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\instruction_reg[3]_i_22_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .I4(\instruction[3]_i_23_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFDF55DFFFDFFFDF))
    \instruction[4]_i_1
       (.I0(\instruction[4]_i_2_n_0 ),
        .I1(\instruction[4]_i_3_n_0 ),
        .I2(\instruction_reg[4]_i_4_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction[4]_i_5_n_0 ),
        .I5(\instruction_reg[4]_i_6_n_0 ),
        .O(\instruction[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAA2AAAAA))
    \instruction[4]_i_12
       (.I0(\instruction_reg[4]_i_25_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\instruction[6]_i_13_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFDFFFFFDFFFFF))
    \instruction[4]_i_14
       (.I0(\instruction[4]_i_28_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[4]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFFDFFFFFFFFDF))
    \instruction[4]_i_15
       (.I0(\instruction[4]_i_29_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[4]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00004498))
    \instruction[4]_i_16
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep_n_0 ),
        .O(\instruction[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h88888888B8888888))
    \instruction[4]_i_17
       (.I0(\instruction_reg[4]_i_30_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\instruction[4]_i_31_n_0 ),
        .I3(\instruction[4]_i_32_n_0 ),
        .I4(\instruction[4]_i_33_n_0 ),
        .I5(\instruction[4]_i_34_n_0 ),
        .O(\instruction[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFD000D0))
    \instruction[4]_i_18
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\instruction[4]_i_35_n_0 ),
        .I2(\instruction_reg[4]_i_36_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[2] ),
        .I4(\instruction[4]_i_37_n_0 ),
        .I5(\instruction[6]_i_31_n_0 ),
        .O(\instruction[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h2210200800800200))
    \instruction[4]_i_19
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000))
    \instruction[4]_i_2
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\instruction[4]_i_7_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[2] ),
        .I3(\instruction[4]_i_8_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\instruction[4]_i_9_n_0 ),
        .O(\instruction[4]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00008244))
    \instruction[4]_i_20
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hF5F7FFF7FFFFFFEF))
    \instruction[4]_i_21
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[4]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF))
    \instruction[4]_i_22
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[4]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFB69BFEFF))
    \instruction[4]_i_23
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[4]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hBBFBBBD9FFF9FBDF))
    \instruction[4]_i_24
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[4]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h28))
    \instruction[4]_i_28
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[4]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[4]_i_29
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h57F7FFFF57F70000))
    \instruction[4]_i_3
       (.I0(\instruction_reg[4]_i_10_n_0 ),
        .I1(\instruction_reg[4]_i_11_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[2] ),
        .I3(\instruction[4]_i_12_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\instruction_reg[4]_i_13_n_0 ),
        .O(\instruction[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFF7FFDFD77D7))
    \instruction[4]_i_31
       (.I0(\instruction[21]_i_30_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDF75DF5F7FF))
    \instruction[4]_i_32
       (.I0(\instruction[25]_i_11_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[4]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7F7F7FFFFFFF))
    \instruction[4]_i_33
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep_n_0_[3] ),
        .I2(\instruction[4]_i_46_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[8] ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000000))
    \instruction[4]_i_34
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[3] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[4]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[4]_i_35
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[4]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA8AAAAAAA))
    \instruction[4]_i_37
       (.I0(\instruction_reg[4]_i_49_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[4]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFDFBF9FFF3DFDFF))
    \instruction[4]_i_38
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hEFEF7EEEFAFFDFFF))
    \instruction[4]_i_39
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[4]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0013050490186004))
    \instruction[4]_i_40
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hA0F00050A0A0548C))
    \instruction[4]_i_41
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[4]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0040051002120210))
    \instruction[4]_i_42
       (.I0(\program_counter_reg_rep_n_0_[2] ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[4]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000000021524200))
    \instruction[4]_i_43
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[4]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFD2FFFFF2FDFF))
    \instruction[4]_i_44
       (.I0(\program_counter_reg_rep_n_0_[3] ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[4]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF6FFF))
    \instruction[4]_i_45
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[3] ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[4]_i_46
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[4]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hF7F7F7F7FBFFFFFB))
    \instruction[4]_i_47
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[4]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFBF7FDAAF6FDEFF5))
    \instruction[4]_i_48
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep_n_0_[8] ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'h20080000))
    \instruction[4]_i_5
       (.I0(\instruction[4]_i_16_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[2] ),
        .O(\instruction[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFD7FFBDFFFDFFD7))
    \instruction[4]_i_50
       (.I0(\program_counter_reg_rep_n_0_[8] ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[4]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEF2FFFF))
    \instruction[4]_i_51
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[4]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000002))
    \instruction[4]_i_7
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[8] ),
        .O(\instruction[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000009000029000))
    \instruction[4]_i_8
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep_n_0_[8] ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF4777FFCF4777))
    \instruction[4]_i_9
       (.I0(\instruction[4]_i_19_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[2] ),
        .I2(\instruction[4]_i_20_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0EFF02FFFFFFFFFF))
    \instruction[5]_i_1
       (.I0(\instruction[5]_i_2_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\instruction[5]_i_3_n_0 ),
        .I4(\instruction_reg[5]_i_4_n_0 ),
        .I5(\instruction_reg[5]_i_5_n_0 ),
        .O(\instruction[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h000000E2E2E200E2))
    \instruction[5]_i_10
       (.I0(\instruction[5]_i_12_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\instruction[5]_i_13_n_0 ),
        .I3(\instruction[5]_i_14_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\instruction_reg[5]_i_15_n_0 ),
        .O(\instruction[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8888AAAAAAAAA))
    \instruction[5]_i_11
       (.I0(\instruction_reg[5]_i_16_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\instruction[2]_i_18_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\instruction[5]_i_17_n_0 ),
        .O(\instruction[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8B888B8B8))
    \instruction[5]_i_12
       (.I0(\instruction_reg[5]_i_18_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction_reg[5]_i_19_n_0 ),
        .I3(\instruction[7]_i_12_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2))
    \instruction[5]_i_13
       (.I0(\instruction[5]_i_20_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\instruction[5]_i_21_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\instruction[5]_i_22_n_0 ),
        .I5(\instruction_reg[5]_i_23_n_0 ),
        .O(\instruction[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0F00000080800000))
    \instruction[5]_i_14
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I3(\instruction[5]_i_24_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0200540400000000))
    \instruction[5]_i_17
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[5]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0800280004000000))
    \instruction[5]_i_2
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I3(\instruction[5]_i_6_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[9] ),
        .I5(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF7FF5FFFF7BEFE))
    \instruction[5]_i_20
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[5]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hEFBFEFE7FFFFEFBF))
    \instruction[5]_i_21
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[5]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFDDBEFFDFDEFEDFB))
    \instruction[5]_i_22
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[5]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h0810))
    \instruction[5]_i_24
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[5]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000284800000000))
    \instruction[5]_i_25
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[5]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000800000000))
    \instruction[5]_i_26
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[5]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA8AAAAA88AAAA))
    \instruction[5]_i_27
       (.I0(\instruction_reg[5]_i_35_n_0 ),
        .I1(\instruction[7]_i_12_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[5]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0000F404F404F404))
    \instruction[5]_i_28
       (.I0(\instruction_reg[5]_i_36_n_0 ),
        .I1(\instruction[5]_i_37_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\instruction_reg[5]_i_38_n_0 ),
        .I4(\instruction[18]_i_34_n_0 ),
        .I5(\instruction[5]_i_39_n_0 ),
        .O(\instruction[5]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBBFE1154FFFFFEF7))
    \instruction[5]_i_29
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[5]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFDFFDFF))
    \instruction[5]_i_3
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\instruction[5]_i_7_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h3CBEFFFBCFEFFCFF))
    \instruction[5]_i_30
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[5]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDBFBD77DA779F))
    \instruction[5]_i_31
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[5]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFF7FFFDFFF7EEF9))
    \instruction[5]_i_32
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[5]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h000000810002A000))
    \instruction[5]_i_33
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .O(\instruction[5]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h8000000001080240))
    \instruction[5]_i_34
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[5]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDFFFFFFEFFFF))
    \instruction[5]_i_37
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[5]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h04))
    \instruction[5]_i_39
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[5]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h88C00300000C4400))
    \instruction[5]_i_42
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[5]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h8889244300006142))
    \instruction[5]_i_43
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[5]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFE65EFFFDEFFEFF))
    \instruction[5]_i_44
       (.I0(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[5]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hF0FDCFFFD3DF13DF))
    \instruction[5]_i_45
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[5]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF7BFC47FFFF))
    \instruction[5]_i_46
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[5]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFBEEFF1))
    \instruction[5]_i_47
       (.I0(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[5]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hBDFBBDFFBDFBBD56))
    \instruction[5]_i_48
       (.I0(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[5]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hEBFEDFEF))
    \instruction[5]_i_49
       (.I0(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[5]_i_49_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[5]_i_6
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFFFBBFFFFFFF))
    \instruction[5]_i_7
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .O(\instruction[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h8C800000B0800008))
    \instruction[5]_i_8
       (.I0(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000))
    \instruction[5]_i_9
       (.I0(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .O(\instruction[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFF8F888FFF8FFF8F))
    \instruction[6]_i_1
       (.I0(\instruction_reg[6]_i_2_n_0 ),
        .I1(\instruction[6]_i_3_n_0 ),
        .I2(\instruction[6]_i_4_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction[6]_i_5_n_0 ),
        .I5(\instruction_reg[6]_i_6_n_0 ),
        .O(\instruction[6]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h9FFF))
    \instruction[6]_i_10
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[6]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h24))
    \instruction[6]_i_12
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[6]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[6]_i_13
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[6]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hE200E2E2E2E2E2E2))
    \instruction[6]_i_14
       (.I0(\instruction[6]_i_26_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\instruction_reg[6]_i_27_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\instruction[6]_i_28_n_0 ),
        .I5(\instruction[6]_i_12_n_0 ),
        .O(\instruction[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFB000B0))
    \instruction[6]_i_15
       (.I0(\instruction[7]_i_12_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\instruction_reg[6]_i_29_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\instruction_reg[6]_i_30_n_0 ),
        .I5(\instruction[6]_i_31_n_0 ),
        .O(\instruction[6]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0009000000000008))
    \instruction[6]_i_16
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .O(\instruction[6]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0090400004001000))
    \instruction[6]_i_17
       (.I0(\program_counter_reg_rep[3]_rep_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000))
    \instruction[6]_i_18
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0028200002808008))
    \instruction[6]_i_19
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[6]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA2AAAA2AAAAA))
    \instruction[6]_i_20
       (.I0(\instruction_reg[6]_i_32_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h800C300080000000))
    \instruction[6]_i_23
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[6]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0040610000000000))
    \instruction[6]_i_24
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[6]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h00000040))
    \instruction[6]_i_25
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hA2AA2AAAAA2AA2AA))
    \instruction[6]_i_26
       (.I0(\instruction_reg[6]_i_37_n_0 ),
        .I1(\instruction[6]_i_13_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[6]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[6]_i_28
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[6]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h6))
    \instruction[6]_i_3
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .O(\instruction[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000224000000000))
    \instruction[6]_i_31
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[3]_rep_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[6]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hEE76BF67F5FFFDEB))
    \instruction[6]_i_33
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[5] ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[6]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hEBE5FBEFFB79FFFD))
    \instruction[6]_i_34
       (.I0(\program_counter_reg_rep_n_0_[5] ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[6]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hEAEEEEEE2A222222))
    \instruction[6]_i_35
       (.I0(\instruction[6]_i_46_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[18]_i_6_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\instruction[6]_i_47_n_0 ),
        .O(\instruction[6]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hE200E2E2E2E2E2E2))
    \instruction[6]_i_36
       (.I0(\instruction[6]_i_48_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[6]_i_49_n_0 ),
        .I3(\instruction[7]_i_12_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hDEFF4E6FFFFD5F7E))
    \instruction[6]_i_38
       (.I0(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[6]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFB4FFFFFCB7FF))
    \instruction[6]_i_39
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[6]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hAA8AA8AAA8AAAAA8))
    \instruction[6]_i_4
       (.I0(\instruction[6]_i_9_n_0 ),
        .I1(\instruction[6]_i_10_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h7D79FD79FFAFDFDF))
    \instruction[6]_i_40
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[6]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFEFEFDEDEFEFD))
    \instruction[6]_i_41
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFF77EE5FEFFEEFFF))
    \instruction[6]_i_42
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[6]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFFFFFFFFFE))
    \instruction[6]_i_43
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[6]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFBCCCFFFFBFFFF))
    \instruction[6]_i_44
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[5] ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[6]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFDBBDFDF2AEF))
    \instruction[6]_i_45
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep_n_0_[5] ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[6]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hDFAADEF56777EFFF))
    \instruction[6]_i_46
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[5] ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[6]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hABFFFFFEFFFFFFBF))
    \instruction[6]_i_47
       (.I0(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFDB9FFFF5F5BFBEB))
    \instruction[6]_i_48
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFDFFFB9E5E5FBFF))
    \instruction[6]_i_49
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h888888888888B888))
    \instruction[6]_i_5
       (.I0(\instruction_reg[6]_i_11_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[6]_i_12_n_0 ),
        .I3(\instruction[6]_i_13_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[5] ),
        .O(\instruction[6]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h722F77FD77F205DF))
    \instruction[6]_i_50
       (.I0(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[6]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFEFFEFEFF))
    \instruction[6]_i_51
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[3]_rep_n_0 ),
        .O(\instruction[6]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFC0))
    \instruction[6]_i_9
       (.I0(\instruction[6]_i_20_n_0 ),
        .I1(\instruction_reg[6]_i_21_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep_n_0 ),
        .I3(\instruction_reg[6]_i_22_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I5(\instruction[6]_i_23_n_0 ),
        .O(\instruction[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7))
    \instruction[7]_i_1
       (.I0(\instruction[7]_i_2_n_0 ),
        .I1(\instruction[7]_i_3_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\instruction[7]_i_4_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\instruction[7]_i_5_n_0 ),
        .O(\instruction[7]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[7]_i_10
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[7]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h80))
    \instruction[7]_i_11
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[7]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[7]_i_12
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[7]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF))
    \instruction[7]_i_13
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[7]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hA1))
    \instruction[7]_i_14
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[7]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h8B8B8BBBBBBB8BBB))
    \instruction[7]_i_16
       (.I0(\instruction[7]_i_23_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\instruction[7]_i_24_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\instruction[7]_i_25_n_0 ),
        .O(\instruction[7]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[7]_i_17
       (.I0(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[7]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFEDEFFFFF5FEF7F))
    \instruction[7]_i_18
       (.I0(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[7]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFBEBBFFFFFFFBFFF))
    \instruction[7]_i_19
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hE7FFFFFFE7FF0000))
    \instruction[7]_i_2
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\instruction[7]_i_6_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\instruction[7]_i_7_n_0 ),
        .O(\instruction[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFDD3FFFFF))
    \instruction[7]_i_20
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .O(\instruction[7]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF))
    \instruction[7]_i_21
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .O(\instruction[7]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAFFBFEFEAFFFFFFF))
    \instruction[7]_i_22
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[7]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h000000001D1D0C3F))
    \instruction[7]_i_23
       (.I0(\instruction[7]_i_26_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\instruction[7]_i_27_n_0 ),
        .I3(\instruction[7]_i_28_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\instruction[7]_i_29_n_0 ),
        .O(\instruction[7]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0000000A00004410))
    \instruction[7]_i_24
       (.I0(\program_counter_reg_rep[2]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[7]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010B80040))
    \instruction[7]_i_25
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .O(\instruction[7]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h4104400400040000))
    \instruction[7]_i_26
       (.I0(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[7]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00A4040000000000))
    \instruction[7]_i_27
       (.I0(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\instruction[7]_i_30_n_0 ),
        .O(\instruction[7]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h8800008000000080))
    \instruction[7]_i_28
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .O(\instruction[7]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000))
    \instruction[7]_i_29
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .O(\instruction[7]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hE2E2E200E2E2E2E2))
    \instruction[7]_i_3
       (.I0(\instruction[7]_i_8_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[1] ),
        .I2(\instruction_reg[7]_i_9_n_0 ),
        .I3(\instruction[7]_i_10_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\instruction[7]_i_11_n_0 ),
        .O(\instruction[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \instruction[7]_i_30
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[7]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hE2FFFFFFE2FF0000))
    \instruction[7]_i_4
       (.I0(\instruction[7]_i_12_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\instruction[7]_i_13_n_0 ),
        .I3(\instruction[7]_i_14_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\instruction_reg[7]_i_15_n_0 ),
        .O(\instruction[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA2AAAAAAA))
    \instruction[7]_i_5
       (.I0(\instruction[7]_i_16_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\program_counter_reg_rep[2]_rep_n_0 ),
        .O(\instruction[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4410000020000000))
    \instruction[7]_i_6
       (.I0(\program_counter_reg_rep_n_0_[4] ),
        .I1(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I5(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .O(\instruction[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFBBFFFFFFFFF))
    \instruction[7]_i_7
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep_n_0 ),
        .I4(\instruction[7]_i_17_n_0 ),
        .I5(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hABFFFFFFABFF0000))
    \instruction[7]_i_8
       (.I0(\instruction[7]_i_17_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep_n_0 ),
        .I5(\instruction[7]_i_18_n_0 ),
        .O(\instruction[7]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB))
    \instruction[8]_i_1
       (.I0(\instruction_reg[8]_i_2_n_0 ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\instruction[8]_i_3_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction[15]_i_5_n_0 ),
        .O(\instruction[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFFBFFFFBFBFF))
    \instruction[8]_i_10
       (.I0(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[8]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBF30B000A0F0A000))
    \instruction[8]_i_11
       (.I0(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[0] ),
        .I2(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2000000))
    \instruction[8]_i_12
       (.I0(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[8]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00004000))
    \instruction[8]_i_13
       (.I0(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hD1F3D1F300F3D1F3))
    \instruction[8]_i_3
       (.I0(\instruction[8]_i_6_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I2(\instruction[15]_i_8_n_0 ),
        .I3(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I5(\instruction[8]_i_7_n_0 ),
        .O(\instruction[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00010000FFFFFFFF))
    \instruction[8]_i_4
       (.I0(\program_counter_reg_rep_n_0_[0] ),
        .I1(\instruction[20]_i_20_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\instruction[8]_i_8_n_0 ),
        .O(\instruction[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h888888B8B8B888B8))
    \instruction[8]_i_5
       (.I0(\instruction_reg[8]_i_9_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[0] ),
        .I2(\instruction[7]_i_14_n_0 ),
        .I3(\instruction[7]_i_12_n_0 ),
        .I4(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .I5(\instruction[7]_i_13_n_0 ),
        .O(\instruction[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAA800A8000804490))
    \instruction[8]_i_6
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .I5(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .O(\instruction[8]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \instruction[8]_i_7
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .O(\instruction[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB800B8FFB8FFB8FF))
    \instruction[8]_i_8
       (.I0(\instruction[15]_i_17_n_0 ),
        .I1(\program_counter_reg_rep_n_0_[0] ),
        .I2(\instruction[8]_i_10_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .I5(\instruction[8]_i_11_n_0 ),
        .O(\instruction[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00008000FFFFFFFF))
    \instruction[9]_i_1
       (.I0(\program_counter_reg_rep[7]_rep_n_0 ),
        .I1(\program_counter_reg_rep[8]_rep_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I4(\instruction[9]_i_2_n_0 ),
        .I5(\instruction[9]_i_3_n_0 ),
        .O(\instruction[9]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h80080008022A0414))
    \instruction[9]_i_10
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[7]_rep_n_0 ),
        .O(\instruction[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h110120210A012021))
    \instruction[9]_i_11
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[7]_rep_n_0 ),
        .I2(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .O(\instruction[9]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBBFFB1E5B1F5))
    \instruction[9]_i_12
       (.I0(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I1(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\program_counter_reg_rep_n_0_[0] ),
        .O(\instruction[9]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h6))
    \instruction[9]_i_13
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[9]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFDBEFFD7))
    \instruction[9]_i_14
       (.I0(\program_counter_reg_rep_n_0_[0] ),
        .I1(\program_counter_reg_rep_n_0_[4] ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I4(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[9]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFB7CBFB))
    \instruction[9]_i_2
       (.I0(\program_counter_reg_rep_n_0_[0] ),
        .I1(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[1] ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .O(\instruction[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h55555555FFFD5555))
    \instruction[9]_i_3
       (.I0(\program_counter_reg_rep[9]_rep_n_0 ),
        .I1(\instruction[9]_i_4_n_0 ),
        .I2(\program_counter_reg_rep[8]_rep_n_0 ),
        .I3(\instruction_reg[9]_i_5_n_0 ),
        .I4(\instruction[9]_i_6_n_0 ),
        .I5(\instruction[9]_i_7_n_0 ),
        .O(\instruction[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA8AAAAAA))
    \instruction[9]_i_4
       (.I0(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[1] ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\program_counter_reg_rep_n_0_[4] ),
        .I5(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .O(\instruction[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hBBBFFFBF))
    \instruction[9]_i_6
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\instruction[9]_i_4_n_0 ),
        .I2(\instruction[9]_i_10_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[0] ),
        .I4(\instruction[9]_i_11_n_0 ),
        .O(\instruction[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00002220AAAA222A))
    \instruction[9]_i_7
       (.I0(\program_counter_reg_rep[8]_rep_n_0 ),
        .I1(\instruction[9]_i_12_n_0 ),
        .I2(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I3(\instruction[9]_i_13_n_0 ),
        .I4(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .I5(\instruction[9]_i_14_n_0 ),
        .O(\instruction[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hD7BEFE3FD7FFEE7F))
    \instruction[9]_i_8
       (.I0(\program_counter_reg_rep_n_0_[1] ),
        .I1(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I3(\program_counter_reg_rep_n_0_[4] ),
        .I4(\program_counter_reg_rep_n_0_[0] ),
        .I5(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .O(\instruction[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hB9ADBE5DED7F177C))
    \instruction[9]_i_9
       (.I0(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .I1(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .I2(\program_counter_reg_rep_n_0_[4] ),
        .I3(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .I4(\program_counter_reg_rep_n_0_[1] ),
        .I5(\program_counter_reg_rep_n_0_[0] ),
        .O(\instruction[9]_i_9_n_0 ));
  FDRE \instruction_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[0]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[0] ),
        .R(1'b0));
  MUXF7 \instruction_reg[0]_i_10
       (.I0(\instruction[0]_i_22_n_0 ),
        .I1(\instruction[0]_i_23_n_0 ),
        .O(\instruction_reg[0]_i_10_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[0]_i_2
       (.I0(\instruction[0]_i_7_n_0 ),
        .I1(\instruction[0]_i_8_n_0 ),
        .O(\instruction_reg[0]_i_2_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[0]_i_20
       (.I0(\instruction[0]_i_41_n_0 ),
        .I1(\instruction[0]_i_42_n_0 ),
        .O(\instruction_reg[0]_i_20_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[0]_i_24
       (.I0(\instruction[0]_i_43_n_0 ),
        .I1(\instruction[0]_i_44_n_0 ),
        .O(\instruction_reg[0]_i_24_n_0 ),
        .S(\program_counter_reg_rep_n_0_[3] ));
  MUXF7 \instruction_reg[0]_i_27
       (.I0(\instruction[0]_i_45_n_0 ),
        .I1(\instruction[0]_i_46_n_0 ),
        .O(\instruction_reg[0]_i_27_n_0 ),
        .S(\program_counter_reg_rep_n_0_[3] ));
  MUXF7 \instruction_reg[0]_i_33
       (.I0(\instruction[0]_i_51_n_0 ),
        .I1(\instruction[0]_i_52_n_0 ),
        .O(\instruction_reg[0]_i_33_n_0 ),
        .S(\program_counter_reg_rep[8]_rep__2_n_0 ));
  MUXF7 \instruction_reg[0]_i_36
       (.I0(\instruction[0]_i_54_n_0 ),
        .I1(\instruction[0]_i_55_n_0 ),
        .O(\instruction_reg[0]_i_36_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[0]_i_37
       (.I0(\instruction[0]_i_56_n_0 ),
        .I1(\instruction[0]_i_57_n_0 ),
        .O(\instruction_reg[0]_i_37_n_0 ),
        .S(\program_counter_reg_rep[8]_rep__1_n_0 ));
  MUXF7 \instruction_reg[0]_i_39
       (.I0(\instruction[0]_i_58_n_0 ),
        .I1(\instruction[0]_i_59_n_0 ),
        .O(\instruction_reg[0]_i_39_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[0]_i_4
       (.I0(\instruction[0]_i_11_n_0 ),
        .I1(\instruction[0]_i_12_n_0 ),
        .O(\instruction_reg[0]_i_4_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[0]_i_47
       (.I0(\instruction[0]_i_60_n_0 ),
        .I1(\instruction[0]_i_61_n_0 ),
        .O(\instruction_reg[0]_i_47_n_0 ),
        .S(\program_counter_reg_rep[7]_rep__0_n_0 ));
  MUXF7 \instruction_reg[0]_i_5
       (.I0(\instruction[0]_i_13_n_0 ),
        .I1(\instruction[0]_i_14_n_0 ),
        .O(\instruction_reg[0]_i_5_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF7 \instruction_reg[0]_i_50
       (.I0(\instruction[0]_i_62_n_0 ),
        .I1(\instruction[0]_i_63_n_0 ),
        .O(\instruction_reg[0]_i_50_n_0 ),
        .S(\program_counter_reg_rep_n_0_[3] ));
  FDRE \instruction_reg[15]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[15]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[15] ),
        .R(1'b0));
  FDRE \instruction_reg[16]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[16]_i_1_n_0 ),
        .Q(address_a[0]),
        .R(1'b0));
  MUXF7 \instruction_reg[16]_i_17
       (.I0(\instruction[16]_i_26_n_0 ),
        .I1(\instruction[16]_i_27_n_0 ),
        .O(\instruction_reg[16]_i_17_n_0 ),
        .S(\program_counter_reg_rep_n_0_[5] ));
  MUXF7 \instruction_reg[16]_i_18
       (.I0(\instruction[16]_i_28_n_0 ),
        .I1(\instruction[16]_i_29_n_0 ),
        .O(\instruction_reg[16]_i_18_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[16]_i_22
       (.I0(\instruction[16]_i_30_n_0 ),
        .I1(\instruction[16]_i_31_n_0 ),
        .O(\instruction_reg[16]_i_22_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[16]_i_3
       (.I0(\instruction[16]_i_8_n_0 ),
        .I1(\instruction[16]_i_9_n_0 ),
        .O(\instruction_reg[16]_i_3_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[16]_i_5
       (.I0(\instruction[16]_i_12_n_0 ),
        .I1(\instruction[16]_i_13_n_0 ),
        .O(\instruction_reg[16]_i_5_n_0 ),
        .S(\program_counter_reg_rep_n_0_[0] ));
  FDRE \instruction_reg[17]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[17]_i_1_n_0 ),
        .Q(address_a[1]),
        .R(1'b0));
  MUXF7 \instruction_reg[17]_i_12
       (.I0(\instruction[17]_i_17_n_0 ),
        .I1(\instruction[17]_i_18_n_0 ),
        .O(\instruction_reg[17]_i_12_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[17]_i_14
       (.I0(\instruction[17]_i_21_n_0 ),
        .I1(\instruction[17]_i_22_n_0 ),
        .O(\instruction_reg[17]_i_14_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[17]_i_26
       (.I0(\instruction[17]_i_42_n_0 ),
        .I1(\instruction[17]_i_43_n_0 ),
        .O(\instruction_reg[17]_i_26_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF7 \instruction_reg[17]_i_3
       (.I0(\instruction[17]_i_8_n_0 ),
        .I1(\instruction[17]_i_9_n_0 ),
        .O(\instruction_reg[17]_i_3_n_0 ),
        .S(\program_counter_reg_rep[7]_rep_n_0 ));
  MUXF7 \instruction_reg[17]_i_30
       (.I0(\instruction[17]_i_44_n_0 ),
        .I1(\instruction[17]_i_45_n_0 ),
        .O(\instruction_reg[17]_i_30_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__1_n_0 ));
  MUXF7 \instruction_reg[17]_i_4
       (.I0(\instruction[17]_i_10_n_0 ),
        .I1(\instruction[17]_i_11_n_0 ),
        .O(\instruction_reg[17]_i_4_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[17]_i_46
       (.I0(\instruction[17]_i_50_n_0 ),
        .I1(\instruction[17]_i_51_n_0 ),
        .O(\instruction_reg[17]_i_46_n_0 ),
        .S(\program_counter_reg_rep[7]_rep_n_0 ));
  FDRE \instruction_reg[18]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[18]_i_1_n_0 ),
        .Q(address_a[2]),
        .R(1'b0));
  MUXF8 \instruction_reg[18]_i_10
       (.I0(\instruction_reg[18]_i_22_n_0 ),
        .I1(\instruction_reg[18]_i_23_n_0 ),
        .O(\instruction_reg[18]_i_10_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[18]_i_12
       (.I0(\instruction[18]_i_27_n_0 ),
        .I1(\instruction[18]_i_28_n_0 ),
        .O(\instruction_reg[18]_i_12_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__1_n_0 ));
  MUXF7 \instruction_reg[18]_i_13
       (.I0(\instruction[18]_i_29_n_0 ),
        .I1(\instruction[18]_i_30_n_0 ),
        .O(\instruction_reg[18]_i_13_n_0 ),
        .S(\program_counter_reg_rep[5]_rep__1_n_0 ));
  MUXF7 \instruction_reg[18]_i_21
       (.I0(\instruction[18]_i_37_n_0 ),
        .I1(\instruction[18]_i_38_n_0 ),
        .O(\instruction_reg[18]_i_21_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[18]_i_22
       (.I0(\instruction[18]_i_39_n_0 ),
        .I1(\instruction[18]_i_40_n_0 ),
        .O(\instruction_reg[18]_i_22_n_0 ),
        .S(\program_counter_reg_rep[9]_rep__2_n_0 ));
  MUXF7 \instruction_reg[18]_i_23
       (.I0(\instruction[18]_i_41_n_0 ),
        .I1(\instruction[18]_i_42_n_0 ),
        .O(\instruction_reg[18]_i_23_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__1_n_0 ));
  MUXF8 \instruction_reg[18]_i_4
       (.I0(\instruction_reg[18]_i_12_n_0 ),
        .I1(\instruction_reg[18]_i_13_n_0 ),
        .O(\instruction_reg[18]_i_4_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[18]_i_5
       (.I0(\instruction[18]_i_14_n_0 ),
        .I1(\instruction[18]_i_15_n_0 ),
        .O(\instruction_reg[18]_i_5_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[18]_i_8
       (.I0(\instruction[18]_i_16_n_0 ),
        .I1(\instruction[18]_i_17_n_0 ),
        .O(\instruction_reg[18]_i_8_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  FDRE \instruction_reg[19]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[19]_i_1_n_0 ),
        .Q(address_a[3]),
        .R(1'b0));
  MUXF7 \instruction_reg[19]_i_10
       (.I0(\instruction[19]_i_19_n_0 ),
        .I1(\instruction[19]_i_20_n_0 ),
        .O(\instruction_reg[19]_i_10_n_0 ),
        .S(\program_counter_reg_rep[6]_rep__0_n_0 ));
  MUXF7 \instruction_reg[19]_i_12
       (.I0(\instruction[19]_i_21_n_0 ),
        .I1(\instruction[19]_i_22_n_0 ),
        .O(\instruction_reg[19]_i_12_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  FDRE \instruction_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[1]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[1] ),
        .R(1'b0));
  MUXF7 \instruction_reg[1]_i_17
       (.I0(\instruction[1]_i_27_n_0 ),
        .I1(\instruction[1]_i_28_n_0 ),
        .O(\instruction_reg[1]_i_17_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[1]_i_18
       (.I0(\instruction[1]_i_29_n_0 ),
        .I1(\instruction[1]_i_30_n_0 ),
        .O(\instruction_reg[1]_i_18_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  MUXF8 \instruction_reg[1]_i_2
       (.I0(\instruction_reg[1]_i_6_n_0 ),
        .I1(\instruction_reg[1]_i_7_n_0 ),
        .O(\instruction_reg[1]_i_2_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[1]_i_23
       (.I0(\instruction[1]_i_42_n_0 ),
        .I1(\instruction[1]_i_43_n_0 ),
        .O(\instruction_reg[1]_i_23_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  MUXF7 \instruction_reg[1]_i_24
       (.I0(\instruction[1]_i_44_n_0 ),
        .I1(\instruction[1]_i_45_n_0 ),
        .O(\instruction_reg[1]_i_24_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[1]_i_4
       (.I0(\instruction[1]_i_8_n_0 ),
        .I1(\instruction[1]_i_9_n_0 ),
        .O(\instruction_reg[1]_i_4_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  MUXF7 \instruction_reg[1]_i_48
       (.I0(\instruction[1]_i_54_n_0 ),
        .I1(\instruction[1]_i_55_n_0 ),
        .O(\instruction_reg[1]_i_48_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  MUXF7 \instruction_reg[1]_i_5
       (.I0(\instruction[1]_i_10_n_0 ),
        .I1(\instruction[1]_i_11_n_0 ),
        .O(\instruction_reg[1]_i_5_n_0 ),
        .S(\program_counter_reg_rep_n_0_[0] ));
  MUXF7 \instruction_reg[1]_i_50
       (.I0(\instruction[1]_i_56_n_0 ),
        .I1(\instruction[1]_i_57_n_0 ),
        .O(\instruction_reg[1]_i_50_n_0 ),
        .S(\program_counter_reg_rep[8]_rep__0_n_0 ));
  MUXF7 \instruction_reg[1]_i_52
       (.I0(\instruction[1]_i_58_n_0 ),
        .I1(\instruction[1]_i_59_n_0 ),
        .O(\instruction_reg[1]_i_52_n_0 ),
        .S(\program_counter_reg_rep_n_0_[6] ));
  MUXF7 \instruction_reg[1]_i_53
       (.I0(\instruction[1]_i_60_n_0 ),
        .I1(\instruction[1]_i_61_n_0 ),
        .O(\instruction_reg[1]_i_53_n_0 ),
        .S(\program_counter_reg_rep[5]_rep__0_n_0 ));
  MUXF7 \instruction_reg[1]_i_6
       (.I0(\instruction[1]_i_12_n_0 ),
        .I1(\instruction[1]_i_13_n_0 ),
        .O(\instruction_reg[1]_i_6_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  MUXF7 \instruction_reg[1]_i_7
       (.I0(\instruction[1]_i_14_n_0 ),
        .I1(\instruction[1]_i_15_n_0 ),
        .O(\instruction_reg[1]_i_7_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  FDRE \instruction_reg[20]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[20]_i_1_n_0 ),
        .Q(address_z[0]),
        .R(1'b0));
  MUXF7 \instruction_reg[20]_i_12
       (.I0(\instruction[20]_i_18_n_0 ),
        .I1(\instruction[20]_i_19_n_0 ),
        .O(\instruction_reg[20]_i_12_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[20]_i_23
       (.I0(\instruction[20]_i_28_n_0 ),
        .I1(\instruction[20]_i_29_n_0 ),
        .O(\instruction_reg[20]_i_23_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF7 \instruction_reg[20]_i_25
       (.I0(\instruction[20]_i_30_n_0 ),
        .I1(\instruction[20]_i_31_n_0 ),
        .O(\instruction_reg[20]_i_25_n_0 ),
        .S(\program_counter_reg_rep_n_0_[3] ));
  MUXF7 \instruction_reg[20]_i_8
       (.I0(\instruction[20]_i_15_n_0 ),
        .I1(\instruction[20]_i_16_n_0 ),
        .O(\instruction_reg[20]_i_8_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  FDRE \instruction_reg[21]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[21]_i_1_n_0 ),
        .Q(address_z[1]),
        .R(1'b0));
  MUXF7 \instruction_reg[21]_i_10
       (.I0(\instruction[21]_i_25_n_0 ),
        .I1(\instruction[21]_i_26_n_0 ),
        .O(\instruction_reg[21]_i_10_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[21]_i_11
       (.I0(\instruction[21]_i_27_n_0 ),
        .I1(\instruction[21]_i_28_n_0 ),
        .O(\instruction_reg[21]_i_11_n_0 ),
        .S(\program_counter_reg_rep_n_0_[3] ));
  MUXF8 \instruction_reg[21]_i_13
       (.I0(\instruction_reg[21]_i_34_n_0 ),
        .I1(\instruction_reg[21]_i_35_n_0 ),
        .O(\instruction_reg[21]_i_13_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__0_n_0 ));
  MUXF7 \instruction_reg[21]_i_33
       (.I0(\instruction[21]_i_47_n_0 ),
        .I1(\instruction[21]_i_48_n_0 ),
        .O(\instruction_reg[21]_i_33_n_0 ),
        .S(\program_counter_reg_rep_n_0_[3] ));
  MUXF7 \instruction_reg[21]_i_34
       (.I0(\instruction[21]_i_49_n_0 ),
        .I1(\instruction[21]_i_50_n_0 ),
        .O(\instruction_reg[21]_i_34_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[21]_i_35
       (.I0(\instruction[21]_i_51_n_0 ),
        .I1(\instruction[21]_i_52_n_0 ),
        .O(\instruction_reg[21]_i_35_n_0 ),
        .S(\program_counter_reg_rep[9]_rep_n_0 ));
  MUXF7 \instruction_reg[21]_i_36
       (.I0(\instruction[21]_i_53_n_0 ),
        .I1(\instruction[21]_i_54_n_0 ),
        .O(\instruction_reg[21]_i_36_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[21]_i_39
       (.I0(\instruction[21]_i_55_n_0 ),
        .I1(\instruction[21]_i_56_n_0 ),
        .O(\instruction_reg[21]_i_39_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[21]_i_4
       (.I0(\instruction[21]_i_14_n_0 ),
        .I1(\instruction[21]_i_15_n_0 ),
        .O(\instruction_reg[21]_i_4_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[21]_i_40
       (.I0(\instruction[21]_i_57_n_0 ),
        .I1(\instruction[21]_i_58_n_0 ),
        .O(\instruction_reg[21]_i_40_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[21]_i_44
       (.I0(\instruction[21]_i_62_n_0 ),
        .I1(\instruction[21]_i_63_n_0 ),
        .O(\instruction_reg[21]_i_44_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[21]_i_5
       (.I0(\instruction[21]_i_16_n_0 ),
        .I1(\instruction[21]_i_17_n_0 ),
        .O(\instruction_reg[21]_i_5_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  FDRE \instruction_reg[22]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[22]_i_1_n_0 ),
        .Q(address_z[2]),
        .R(1'b0));
  MUXF7 \instruction_reg[22]_i_5
       (.I0(\instruction[22]_i_9_n_0 ),
        .I1(\instruction[22]_i_10_n_0 ),
        .O(\instruction_reg[22]_i_5_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  FDRE \instruction_reg[23]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[23]_i_1_n_0 ),
        .Q(address_z[3]),
        .R(1'b0));
  MUXF7 \instruction_reg[23]_i_10
       (.I0(\instruction[23]_i_20_n_0 ),
        .I1(\instruction[23]_i_21_n_0 ),
        .O(\instruction_reg[23]_i_10_n_0 ),
        .S(\program_counter_reg_rep[6]_rep__0_n_0 ));
  MUXF7 \instruction_reg[23]_i_2
       (.I0(\instruction[23]_i_7_n_0 ),
        .I1(\instruction[23]_i_8_n_0 ),
        .O(\instruction_reg[23]_i_2_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF8 \instruction_reg[23]_i_27
       (.I0(\instruction_reg[23]_i_44_n_0 ),
        .I1(\instruction_reg[23]_i_45_n_0 ),
        .O(\instruction_reg[23]_i_27_n_0 ),
        .S(\program_counter_reg_rep[9]_rep__1_n_0 ));
  MUXF7 \instruction_reg[23]_i_33
       (.I0(\instruction[23]_i_48_n_0 ),
        .I1(\instruction[23]_i_49_n_0 ),
        .O(\instruction_reg[23]_i_33_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[23]_i_4
       (.I0(\instruction[23]_i_12_n_0 ),
        .I1(\instruction[23]_i_13_n_0 ),
        .O(\instruction_reg[23]_i_4_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[23]_i_40
       (.I0(\instruction[23]_i_50_n_0 ),
        .I1(\instruction[23]_i_51_n_0 ),
        .O(\instruction_reg[23]_i_40_n_0 ),
        .S(\program_counter_reg_rep[9]_rep__1_n_0 ));
  MUXF7 \instruction_reg[23]_i_43
       (.I0(\instruction[23]_i_52_n_0 ),
        .I1(\instruction[23]_i_53_n_0 ),
        .O(\instruction_reg[23]_i_43_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[23]_i_44
       (.I0(\instruction[23]_i_54_n_0 ),
        .I1(\instruction[23]_i_55_n_0 ),
        .O(\instruction_reg[23]_i_44_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF7 \instruction_reg[23]_i_45
       (.I0(\instruction[23]_i_56_n_0 ),
        .I1(\instruction[23]_i_57_n_0 ),
        .O(\instruction_reg[23]_i_45_n_0 ),
        .S(\program_counter_reg_rep[5]_rep_n_0 ));
  MUXF7 \instruction_reg[23]_i_5
       (.I0(\instruction[23]_i_14_n_0 ),
        .I1(\instruction[23]_i_15_n_0 ),
        .O(\instruction_reg[23]_i_5_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[23]_i_6
       (.I0(\instruction[23]_i_16_n_0 ),
        .I1(\instruction[23]_i_17_n_0 ),
        .O(\instruction_reg[23]_i_6_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  FDRE \instruction_reg[24]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[24]_i_1_n_0 ),
        .Q(opcode[0]),
        .R(1'b0));
  MUXF7 \instruction_reg[24]_i_19
       (.I0(\instruction[24]_i_34_n_0 ),
        .I1(\instruction[24]_i_35_n_0 ),
        .O(\instruction_reg[24]_i_19_n_0 ),
        .S(\program_counter_reg_rep[9]_rep_n_0 ));
  MUXF7 \instruction_reg[24]_i_20
       (.I0(\instruction[24]_i_36_n_0 ),
        .I1(\instruction[24]_i_37_n_0 ),
        .O(\instruction_reg[24]_i_20_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[24]_i_25
       (.I0(\instruction[24]_i_47_n_0 ),
        .I1(\instruction[24]_i_48_n_0 ),
        .O(\instruction_reg[24]_i_25_n_0 ),
        .S(\program_counter_reg_rep[5]_rep__2_n_0 ));
  MUXF7 \instruction_reg[24]_i_3
       (.I0(\instruction[24]_i_7_n_0 ),
        .I1(\instruction[24]_i_8_n_0 ),
        .O(\instruction_reg[24]_i_3_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[24]_i_4
       (.I0(\instruction[24]_i_9_n_0 ),
        .I1(\instruction[24]_i_10_n_0 ),
        .O(\instruction_reg[24]_i_4_n_0 ),
        .S(\program_counter_reg_rep[8]_rep_n_0 ));
  MUXF7 \instruction_reg[24]_i_41
       (.I0(\instruction[24]_i_53_n_0 ),
        .I1(\instruction[24]_i_54_n_0 ),
        .O(\instruction_reg[24]_i_41_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[24]_i_45
       (.I0(\instruction[24]_i_55_n_0 ),
        .I1(\instruction[24]_i_56_n_0 ),
        .O(\instruction_reg[24]_i_45_n_0 ),
        .S(\program_counter_reg_rep_n_0_[6] ));
  MUXF7 \instruction_reg[24]_i_5
       (.I0(\instruction[24]_i_11_n_0 ),
        .I1(\instruction[24]_i_12_n_0 ),
        .O(\instruction_reg[24]_i_5_n_0 ),
        .S(\program_counter_reg_rep_n_0_[0] ));
  FDRE \instruction_reg[25]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[25]_i_1_n_0 ),
        .Q(opcode[1]),
        .R(1'b0));
  MUXF8 \instruction_reg[25]_i_19
       (.I0(\instruction_reg[25]_i_31_n_0 ),
        .I1(\instruction_reg[25]_i_32_n_0 ),
        .O(\instruction_reg[25]_i_19_n_0 ),
        .S(\instruction[25]_i_30_n_0 ));
  MUXF8 \instruction_reg[25]_i_20
       (.I0(\instruction_reg[25]_i_33_n_0 ),
        .I1(\instruction_reg[25]_i_34_n_0 ),
        .O(\instruction_reg[25]_i_20_n_0 ),
        .S(\program_counter_reg_rep[9]_rep__1_n_0 ));
  MUXF7 \instruction_reg[25]_i_26
       (.I0(\instruction[25]_i_36_n_0 ),
        .I1(\instruction[25]_i_37_n_0 ),
        .O(\instruction_reg[25]_i_26_n_0 ),
        .S(\program_counter_reg_rep_n_0_[7] ));
  MUXF7 \instruction_reg[25]_i_31
       (.I0(\instruction[25]_i_40_n_0 ),
        .I1(\instruction[25]_i_41_n_0 ),
        .O(\instruction_reg[25]_i_31_n_0 ),
        .S(\program_counter_reg_rep[4]_rep_n_0 ));
  MUXF7 \instruction_reg[25]_i_32
       (.I0(\instruction[25]_i_42_n_0 ),
        .I1(\instruction[25]_i_43_n_0 ),
        .O(\instruction_reg[25]_i_32_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[25]_i_33
       (.I0(\instruction[25]_i_44_n_0 ),
        .I1(\instruction[25]_i_45_n_0 ),
        .O(\instruction_reg[25]_i_33_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[25]_i_34
       (.I0(\instruction[25]_i_46_n_0 ),
        .I1(\instruction[25]_i_47_n_0 ),
        .O(\instruction_reg[25]_i_34_n_0 ),
        .S(\program_counter_reg_rep_n_0_[3] ));
  MUXF7 \instruction_reg[25]_i_4
       (.I0(\instruction[25]_i_12_n_0 ),
        .I1(\instruction[25]_i_13_n_0 ),
        .O(\instruction_reg[25]_i_4_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  FDRE \instruction_reg[26]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[26]_i_1_n_0 ),
        .Q(opcode[2]),
        .R(1'b0));
  MUXF7 \instruction_reg[26]_i_10
       (.I0(\instruction[26]_i_15_n_0 ),
        .I1(\instruction[26]_i_16_n_0 ),
        .O(\instruction_reg[26]_i_10_n_0 ),
        .S(\program_counter_reg_rep_n_0_[7] ));
  MUXF7 \instruction_reg[26]_i_21
       (.I0(\instruction[26]_i_24_n_0 ),
        .I1(\instruction[26]_i_25_n_0 ),
        .O(\instruction_reg[26]_i_21_n_0 ),
        .S(\program_counter_reg_rep_n_0_[4] ));
  FDRE \instruction_reg[27]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[27]_i_1_n_0 ),
        .Q(opcode[3]),
        .R(1'b0));
  MUXF7 \instruction_reg[27]_i_12
       (.I0(\instruction[27]_i_14_n_0 ),
        .I1(\instruction[27]_i_15_n_0 ),
        .O(\instruction_reg[27]_i_12_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[27]_i_3
       (.I0(\instruction[27]_i_4_n_0 ),
        .I1(\instruction[27]_i_5_n_0 ),
        .O(\instruction_reg[27]_i_3_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  FDRE \instruction_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[2]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[2] ),
        .R(1'b0));
  MUXF7 \instruction_reg[2]_i_16
       (.I0(\instruction[2]_i_34_n_0 ),
        .I1(\instruction[2]_i_35_n_0 ),
        .O(\instruction_reg[2]_i_16_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF8 \instruction_reg[2]_i_19
       (.I0(\instruction_reg[2]_i_37_n_0 ),
        .I1(\instruction_reg[2]_i_38_n_0 ),
        .O(\instruction_reg[2]_i_19_n_0 ),
        .S(\instruction[2]_i_36_n_0 ));
  MUXF7 \instruction_reg[2]_i_2
       (.I0(\instruction[2]_i_7_n_0 ),
        .I1(\instruction[2]_i_8_n_0 ),
        .O(\instruction_reg[2]_i_2_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[2]_i_28
       (.I0(\instruction[2]_i_41_n_0 ),
        .I1(\instruction[2]_i_42_n_0 ),
        .O(\instruction_reg[2]_i_28_n_0 ),
        .S(\program_counter_reg_rep[9]_rep__0_n_0 ));
  MUXF7 \instruction_reg[2]_i_30
       (.I0(\instruction[2]_i_43_n_0 ),
        .I1(\instruction[2]_i_44_n_0 ),
        .O(\instruction_reg[2]_i_30_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__0_n_0 ));
  MUXF7 \instruction_reg[2]_i_31
       (.I0(\instruction[2]_i_45_n_0 ),
        .I1(\instruction[2]_i_46_n_0 ),
        .O(\instruction_reg[2]_i_31_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__0_n_0 ));
  MUXF7 \instruction_reg[2]_i_37
       (.I0(\instruction[2]_i_51_n_0 ),
        .I1(\instruction[2]_i_52_n_0 ),
        .O(\instruction_reg[2]_i_37_n_0 ),
        .S(\program_counter_reg_rep[7]_rep__1_n_0 ));
  MUXF7 \instruction_reg[2]_i_38
       (.I0(\instruction[2]_i_53_n_0 ),
        .I1(\instruction[2]_i_54_n_0 ),
        .O(\instruction_reg[2]_i_38_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__1_n_0 ));
  MUXF7 \instruction_reg[2]_i_4
       (.I0(\instruction[2]_i_12_n_0 ),
        .I1(\instruction[2]_i_13_n_0 ),
        .O(\instruction_reg[2]_i_4_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[2]_i_48
       (.I0(\instruction[2]_i_55_n_0 ),
        .I1(\instruction[2]_i_56_n_0 ),
        .O(\instruction_reg[2]_i_48_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__0_n_0 ));
  MUXF7 \instruction_reg[2]_i_5
       (.I0(\instruction[2]_i_14_n_0 ),
        .I1(\instruction[2]_i_15_n_0 ),
        .O(\instruction_reg[2]_i_5_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  FDRE \instruction_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[3]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[3] ),
        .R(1'b0));
  MUXF7 \instruction_reg[3]_i_13
       (.I0(\instruction[3]_i_25_n_0 ),
        .I1(\instruction[3]_i_26_n_0 ),
        .O(\instruction_reg[3]_i_13_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[3]_i_14
       (.I0(\instruction[3]_i_27_n_0 ),
        .I1(\instruction[3]_i_28_n_0 ),
        .O(\instruction_reg[3]_i_14_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF7 \instruction_reg[3]_i_17
       (.I0(\instruction[3]_i_37_n_0 ),
        .I1(\instruction[3]_i_38_n_0 ),
        .O(\instruction_reg[3]_i_17_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[3]_i_18
       (.I0(\instruction[3]_i_39_n_0 ),
        .I1(\instruction[3]_i_40_n_0 ),
        .O(\instruction_reg[3]_i_18_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__2_n_0 ));
  MUXF7 \instruction_reg[3]_i_22
       (.I0(\instruction[3]_i_42_n_0 ),
        .I1(\instruction[3]_i_43_n_0 ),
        .O(\instruction_reg[3]_i_22_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF7 \instruction_reg[3]_i_24
       (.I0(\instruction[3]_i_44_n_0 ),
        .I1(\instruction[3]_i_45_n_0 ),
        .O(\instruction_reg[3]_i_24_n_0 ),
        .S(\program_counter_reg_rep_n_0_[6] ));
  MUXF7 \instruction_reg[3]_i_3
       (.I0(\instruction[3]_i_9_n_0 ),
        .I1(\instruction[3]_i_10_n_0 ),
        .O(\instruction_reg[3]_i_3_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[3]_i_5
       (.I0(\instruction[3]_i_15_n_0 ),
        .I1(\instruction[3]_i_16_n_0 ),
        .O(\instruction_reg[3]_i_5_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[3]_i_52
       (.I0(\instruction[3]_i_69_n_0 ),
        .I1(\instruction[3]_i_70_n_0 ),
        .O(\instruction_reg[3]_i_52_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[3]_i_53
       (.I0(\instruction[3]_i_71_n_0 ),
        .I1(\instruction[3]_i_72_n_0 ),
        .O(\instruction_reg[3]_i_53_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__2_n_0 ));
  MUXF7 \instruction_reg[3]_i_56
       (.I0(\instruction[3]_i_76_n_0 ),
        .I1(\instruction[3]_i_77_n_0 ),
        .O(\instruction_reg[3]_i_56_n_0 ),
        .S(\program_counter_reg_rep[8]_rep__0_n_0 ));
  MUXF7 \instruction_reg[3]_i_57
       (.I0(\instruction[3]_i_78_n_0 ),
        .I1(\instruction[3]_i_79_n_0 ),
        .O(\instruction_reg[3]_i_57_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF7 \instruction_reg[3]_i_59
       (.I0(\instruction[3]_i_80_n_0 ),
        .I1(\instruction[3]_i_81_n_0 ),
        .O(\instruction_reg[3]_i_59_n_0 ),
        .S(\program_counter_reg_rep[2]_rep_n_0 ));
  MUXF7 \instruction_reg[3]_i_65
       (.I0(\instruction[3]_i_82_n_0 ),
        .I1(\instruction[3]_i_83_n_0 ),
        .O(\instruction_reg[3]_i_65_n_0 ),
        .S(\program_counter_reg_rep[7]_rep__1_n_0 ));
  FDRE \instruction_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[4]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[4] ),
        .R(1'b0));
  MUXF7 \instruction_reg[4]_i_10
       (.I0(\instruction[4]_i_21_n_0 ),
        .I1(\instruction[4]_i_22_n_0 ),
        .O(\instruction_reg[4]_i_10_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[4]_i_11
       (.I0(\instruction[4]_i_23_n_0 ),
        .I1(\instruction[4]_i_24_n_0 ),
        .O(\instruction_reg[4]_i_11_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF8 \instruction_reg[4]_i_13
       (.I0(\instruction_reg[4]_i_26_n_0 ),
        .I1(\instruction_reg[4]_i_27_n_0 ),
        .O(\instruction_reg[4]_i_13_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[4]_i_25
       (.I0(\instruction[4]_i_38_n_0 ),
        .I1(\instruction[4]_i_39_n_0 ),
        .O(\instruction_reg[4]_i_25_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[4]_i_26
       (.I0(\instruction[4]_i_40_n_0 ),
        .I1(\instruction[4]_i_41_n_0 ),
        .O(\instruction_reg[4]_i_26_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[4]_i_27
       (.I0(\instruction[4]_i_42_n_0 ),
        .I1(\instruction[4]_i_43_n_0 ),
        .O(\instruction_reg[4]_i_27_n_0 ),
        .S(\program_counter_reg_rep[7]_rep__0_n_0 ));
  MUXF7 \instruction_reg[4]_i_30
       (.I0(\instruction[4]_i_44_n_0 ),
        .I1(\instruction[4]_i_45_n_0 ),
        .O(\instruction_reg[4]_i_30_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[4]_i_36
       (.I0(\instruction[4]_i_47_n_0 ),
        .I1(\instruction[4]_i_48_n_0 ),
        .O(\instruction_reg[4]_i_36_n_0 ),
        .S(\program_counter_reg_rep_n_0_[4] ));
  MUXF7 \instruction_reg[4]_i_4
       (.I0(\instruction[4]_i_14_n_0 ),
        .I1(\instruction[4]_i_15_n_0 ),
        .O(\instruction_reg[4]_i_4_n_0 ),
        .S(\program_counter_reg_rep_n_0_[2] ));
  MUXF7 \instruction_reg[4]_i_49
       (.I0(\instruction[4]_i_50_n_0 ),
        .I1(\instruction[4]_i_51_n_0 ),
        .O(\instruction_reg[4]_i_49_n_0 ),
        .S(\program_counter_reg_rep_n_0_[4] ));
  MUXF7 \instruction_reg[4]_i_6
       (.I0(\instruction[4]_i_17_n_0 ),
        .I1(\instruction[4]_i_18_n_0 ),
        .O(\instruction_reg[4]_i_6_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  FDRE \instruction_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[5]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[5] ),
        .R(1'b0));
  MUXF7 \instruction_reg[5]_i_15
       (.I0(\instruction[5]_i_25_n_0 ),
        .I1(\instruction[5]_i_26_n_0 ),
        .O(\instruction_reg[5]_i_15_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__0_n_0 ));
  MUXF7 \instruction_reg[5]_i_16
       (.I0(\instruction[5]_i_27_n_0 ),
        .I1(\instruction[5]_i_28_n_0 ),
        .O(\instruction_reg[5]_i_16_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[5]_i_18
       (.I0(\instruction[5]_i_29_n_0 ),
        .I1(\instruction[5]_i_30_n_0 ),
        .O(\instruction_reg[5]_i_18_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__0_n_0 ));
  MUXF7 \instruction_reg[5]_i_19
       (.I0(\instruction[5]_i_31_n_0 ),
        .I1(\instruction[5]_i_32_n_0 ),
        .O(\instruction_reg[5]_i_19_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__1_n_0 ));
  MUXF7 \instruction_reg[5]_i_23
       (.I0(\instruction[5]_i_33_n_0 ),
        .I1(\instruction[5]_i_34_n_0 ),
        .O(\instruction_reg[5]_i_23_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF8 \instruction_reg[5]_i_35
       (.I0(\instruction_reg[5]_i_40_n_0 ),
        .I1(\instruction_reg[5]_i_41_n_0 ),
        .O(\instruction_reg[5]_i_35_n_0 ),
        .S(\program_counter_reg_rep[7]_rep__0_n_0 ));
  MUXF7 \instruction_reg[5]_i_36
       (.I0(\instruction[5]_i_42_n_0 ),
        .I1(\instruction[5]_i_43_n_0 ),
        .O(\instruction_reg[5]_i_36_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__0_n_0 ));
  MUXF7 \instruction_reg[5]_i_38
       (.I0(\instruction[5]_i_44_n_0 ),
        .I1(\instruction[5]_i_45_n_0 ),
        .O(\instruction_reg[5]_i_38_n_0 ),
        .S(\program_counter_reg_rep[7]_rep__0_n_0 ));
  MUXF7 \instruction_reg[5]_i_4
       (.I0(\instruction[5]_i_8_n_0 ),
        .I1(\instruction[5]_i_9_n_0 ),
        .O(\instruction_reg[5]_i_4_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__0_n_0 ));
  MUXF7 \instruction_reg[5]_i_40
       (.I0(\instruction[5]_i_46_n_0 ),
        .I1(\instruction[5]_i_47_n_0 ),
        .O(\instruction_reg[5]_i_40_n_0 ),
        .S(\program_counter_reg_rep[4]_rep__1_n_0 ));
  MUXF7 \instruction_reg[5]_i_41
       (.I0(\instruction[5]_i_48_n_0 ),
        .I1(\instruction[5]_i_49_n_0 ),
        .O(\instruction_reg[5]_i_41_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__0_n_0 ));
  MUXF7 \instruction_reg[5]_i_5
       (.I0(\instruction[5]_i_10_n_0 ),
        .I1(\instruction[5]_i_11_n_0 ),
        .O(\instruction_reg[5]_i_5_n_0 ),
        .S(\program_counter_reg_rep_n_0_[0] ));
  FDRE \instruction_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[6]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[6] ),
        .R(1'b0));
  MUXF7 \instruction_reg[6]_i_11
       (.I0(\instruction[6]_i_24_n_0 ),
        .I1(\instruction[6]_i_25_n_0 ),
        .O(\instruction_reg[6]_i_11_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF8 \instruction_reg[6]_i_2
       (.I0(\instruction_reg[6]_i_7_n_0 ),
        .I1(\instruction_reg[6]_i_8_n_0 ),
        .O(\instruction_reg[6]_i_2_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[6]_i_21
       (.I0(\instruction[6]_i_33_n_0 ),
        .I1(\instruction[6]_i_34_n_0 ),
        .O(\instruction_reg[6]_i_21_n_0 ),
        .S(\program_counter_reg_rep[7]_rep__0_n_0 ));
  MUXF7 \instruction_reg[6]_i_22
       (.I0(\instruction[6]_i_35_n_0 ),
        .I1(\instruction[6]_i_36_n_0 ),
        .O(\instruction_reg[6]_i_22_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[6]_i_27
       (.I0(\instruction[6]_i_38_n_0 ),
        .I1(\instruction[6]_i_39_n_0 ),
        .O(\instruction_reg[6]_i_27_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[6]_i_29
       (.I0(\instruction[6]_i_40_n_0 ),
        .I1(\instruction[6]_i_41_n_0 ),
        .O(\instruction_reg[6]_i_29_n_0 ),
        .S(\program_counter_reg_rep[3]_rep_n_0 ));
  MUXF7 \instruction_reg[6]_i_30
       (.I0(\instruction[6]_i_42_n_0 ),
        .I1(\instruction[6]_i_43_n_0 ),
        .O(\instruction_reg[6]_i_30_n_0 ),
        .S(\program_counter_reg_rep_n_0_[5] ));
  MUXF7 \instruction_reg[6]_i_32
       (.I0(\instruction[6]_i_44_n_0 ),
        .I1(\instruction[6]_i_45_n_0 ),
        .O(\instruction_reg[6]_i_32_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[6]_i_37
       (.I0(\instruction[6]_i_50_n_0 ),
        .I1(\instruction[6]_i_51_n_0 ),
        .O(\instruction_reg[6]_i_37_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[6]_i_6
       (.I0(\instruction[6]_i_14_n_0 ),
        .I1(\instruction[6]_i_15_n_0 ),
        .O(\instruction_reg[6]_i_6_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  MUXF7 \instruction_reg[6]_i_7
       (.I0(\instruction[6]_i_16_n_0 ),
        .I1(\instruction[6]_i_17_n_0 ),
        .O(\instruction_reg[6]_i_7_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  MUXF7 \instruction_reg[6]_i_8
       (.I0(\instruction[6]_i_18_n_0 ),
        .I1(\instruction[6]_i_19_n_0 ),
        .O(\instruction_reg[6]_i_8_n_0 ),
        .S(\program_counter_reg_rep[2]_rep__0_n_0 ));
  FDRE \instruction_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[7]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[7] ),
        .R(1'b0));
  MUXF7 \instruction_reg[7]_i_15
       (.I0(\instruction[7]_i_21_n_0 ),
        .I1(\instruction[7]_i_22_n_0 ),
        .O(\instruction_reg[7]_i_15_n_0 ),
        .S(\program_counter_reg_rep[6]_rep__2_n_0 ));
  MUXF7 \instruction_reg[7]_i_9
       (.I0(\instruction[7]_i_19_n_0 ),
        .I1(\instruction[7]_i_20_n_0 ),
        .O(\instruction_reg[7]_i_9_n_0 ),
        .S(\program_counter_reg_rep_n_0_[4] ));
  FDRE \instruction_reg[8]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[8]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[8] ),
        .R(1'b0));
  MUXF7 \instruction_reg[8]_i_2
       (.I0(\instruction[8]_i_4_n_0 ),
        .I1(\instruction[8]_i_5_n_0 ),
        .O(\instruction_reg[8]_i_2_n_0 ),
        .S(\program_counter_reg_rep[3]_rep__1_n_0 ));
  MUXF7 \instruction_reg[8]_i_9
       (.I0(\instruction[8]_i_12_n_0 ),
        .I1(\instruction[8]_i_13_n_0 ),
        .O(\instruction_reg[8]_i_9_n_0 ),
        .S(\program_counter_reg_rep_n_0_[1] ));
  FDRE \instruction_reg[9]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\instruction[9]_i_1_n_0 ),
        .Q(\instruction_reg_n_0_[9] ),
        .R(1'b0));
  MUXF7 \instruction_reg[9]_i_5
       (.I0(\instruction[9]_i_8_n_0 ),
        .I1(\instruction[9]_i_9_n_0 ),
        .O(\instruction_reg[9]_i_5_n_0 ),
        .S(\program_counter_reg_rep[7]_rep_n_0 ));
  FDRE \literal_2_reg[15]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[15] ),
        .Q(literal_2[15]),
        .R(1'b0));
  FDRE \literal_2_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[4] ),
        .Q(literal_2[4]),
        .R(1'b0));
  FDRE \literal_2_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[5] ),
        .Q(literal_2[5]),
        .R(1'b0));
  FDRE \literal_2_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[6] ),
        .Q(literal_2[6]),
        .R(1'b0));
  FDRE \literal_2_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[7] ),
        .Q(literal_2[7]),
        .R(1'b0));
  FDRE \literal_2_reg[8]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[8] ),
        .Q(literal_2[8]),
        .R(1'b0));
  FDRE \literal_2_reg[9]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(\instruction_reg_n_0_[9] ),
        .Q(literal_2[9]),
        .R(1'b0));
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *)
  (* RTL_RAM_BITS = "131104" *)
  (* RTL_RAM_NAME = "memory" *)
  (* bram_addr_begin = "0" *)
  (* bram_addr_end = "8191" *)
  (* bram_slice_begin = "0" *)
  (* bram_slice_end = "3" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(0))
    memory_reg_0
       (.ADDRARDADDR({1'b1,\write_output[12]_i_1_n_0 ,\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 ,\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 ,\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 ,1'b1,1'b1}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .CASCADEINA(1'b1),
        .CASCADEINB(1'b0),
        .CASCADEOUTA(NLW_memory_reg_0_CASCADEOUTA_UNCONNECTED),
        .CASCADEOUTB(NLW_memory_reg_0_CASCADEOUTB_UNCONNECTED),
        .CLKARDCLK(ETH_CLK_OBUF),
        .CLKBWRCLK(1'b0),
        .DBITERR(NLW_memory_reg_0_DBITERR_UNCONNECTED),
        .DIADI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,store_data[3:0]}),
        .DIBDI({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DIPADIP({1'b0,1'b0,1'b0,1'b0}),
        .DIPBDIP({1'b1,1'b1,1'b1,1'b1}),
        .DOADO({NLW_memory_reg_0_DOADO_UNCONNECTED[31:4],load_data[3:0]}),
        .DOBDO(NLW_memory_reg_0_DOBDO_UNCONNECTED[31:0]),
        .DOPADOP(NLW_memory_reg_0_DOPADOP_UNCONNECTED[3:0]),
        .DOPBDOP(NLW_memory_reg_0_DOPBDOP_UNCONNECTED[3:0]),
        .ECCPARITY(NLW_memory_reg_0_ECCPARITY_UNCONNECTED[7:0]),
        .ENARDEN(1'b1),
        .ENBWREN(1'b0),
        .INJECTDBITERR(NLW_memory_reg_0_INJECTDBITERR_UNCONNECTED),
        .INJECTSBITERR(NLW_memory_reg_0_INJECTSBITERR_UNCONNECTED),
        .RDADDRECC(NLW_memory_reg_0_RDADDRECC_UNCONNECTED[8:0]),
        .REGCEAREGCE(NLW_memory_reg_0_REGCEAREGCE_UNCONNECTED),
        .REGCEB(NLW_memory_reg_0_REGCEB_UNCONNECTED),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SBITERR(NLW_memory_reg_0_SBITERR_UNCONNECTED),
        .WEA({1'b0,1'b0,1'b0,p_0_in}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
  LUT5 #(
    .INIT(32'h00400000))
    memory_reg_0_i_1
       (.I0(\state_reg_n_0_[2] ),
        .I1(\state_reg_n_0_[1] ),
        .I2(opcode_2[1]),
        .I3(opcode_2[0]),
        .I4(memory_reg_0_i_2_n_0),
        .O(p_0_in));
  LUT3 #(
    .INIT(8'h04))
    memory_reg_0_i_2
       (.I0(opcode_2[2]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[3]),
        .O(memory_reg_0_i_2_n_0));
  (* IS_CLOCK_GATED *)
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *)
  (* POWER_OPTED_CE = "ENARDEN=NEW" *)
  (* RTL_RAM_BITS = "131104" *)
  (* RTL_RAM_NAME = "memory" *)
  (* bram_addr_begin = "0" *)
  (* bram_addr_end = "8191" *)
  (* bram_slice_begin = "4" *)
  (* bram_slice_end = "7" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(0))
    memory_reg_1
       (.ADDRARDADDR({1'b1,\write_output[12]_i_1_n_0 ,\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 ,\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 ,\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 ,1'b1,1'b1}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .CASCADEINA(1'b1),
        .CASCADEINB(1'b0),
        .CASCADEOUTA(NLW_memory_reg_1_CASCADEOUTA_UNCONNECTED),
        .CASCADEOUTB(NLW_memory_reg_1_CASCADEOUTB_UNCONNECTED),
        .CLKARDCLK(ETH_CLK_OBUF),
        .CLKBWRCLK(1'b0),
        .DBITERR(NLW_memory_reg_1_DBITERR_UNCONNECTED),
        .DIADI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,store_data[7:4]}),
        .DIBDI({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DIPADIP({1'b0,1'b0,1'b0,1'b0}),
        .DIPBDIP({1'b1,1'b1,1'b1,1'b1}),
        .DOADO({NLW_memory_reg_1_DOADO_UNCONNECTED[31:4],load_data[7:4]}),
        .DOBDO(NLW_memory_reg_1_DOBDO_UNCONNECTED[31:0]),
        .DOPADOP(NLW_memory_reg_1_DOPADOP_UNCONNECTED[3:0]),
        .DOPBDOP(NLW_memory_reg_1_DOPBDOP_UNCONNECTED[3:0]),
        .ECCPARITY(NLW_memory_reg_1_ECCPARITY_UNCONNECTED[7:0]),
        .ENARDEN(memory_reg_1_ENARDEN_cooolgate_en_sig_1),
        .ENBWREN(1'b0),
        .INJECTDBITERR(NLW_memory_reg_1_INJECTDBITERR_UNCONNECTED),
        .INJECTSBITERR(NLW_memory_reg_1_INJECTSBITERR_UNCONNECTED),
        .RDADDRECC(NLW_memory_reg_1_RDADDRECC_UNCONNECTED[8:0]),
        .REGCEAREGCE(NLW_memory_reg_1_REGCEAREGCE_UNCONNECTED),
        .REGCEB(NLW_memory_reg_1_REGCEB_UNCONNECTED),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SBITERR(NLW_memory_reg_1_SBITERR_UNCONNECTED),
        .WEA({1'b0,1'b0,1'b0,p_0_in}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
  LUT4 #(
    .INIT(16'hff02))
    memory_reg_1_ENARDEN_cooolgate_en_gate_1
       (.I0(\state[2]_i_1_n_0 ),
        .I1(\state[0]_i_1_n_0 ),
        .I2(INTERNAL_RST_reg),
        .I3(p_0_in),
        .O(memory_reg_1_ENARDEN_cooolgate_en_sig_1));
  (* IS_CLOCK_GATED *)
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *)
  (* POWER_OPTED_CE = "ENARDEN=NEW" *)
  (* RTL_RAM_BITS = "131104" *)
  (* RTL_RAM_NAME = "memory" *)
  (* bram_addr_begin = "0" *)
  (* bram_addr_end = "8191" *)
  (* bram_slice_begin = "8" *)
  (* bram_slice_end = "11" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(0))
    memory_reg_2
       (.ADDRARDADDR({1'b1,\write_output[12]_i_1_n_0 ,\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 ,\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 ,\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 ,1'b1,1'b1}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .CASCADEINA(1'b1),
        .CASCADEINB(1'b0),
        .CASCADEOUTA(NLW_memory_reg_2_CASCADEOUTA_UNCONNECTED),
        .CASCADEOUTB(NLW_memory_reg_2_CASCADEOUTB_UNCONNECTED),
        .CLKARDCLK(ETH_CLK_OBUF),
        .CLKBWRCLK(1'b0),
        .DBITERR(NLW_memory_reg_2_DBITERR_UNCONNECTED),
        .DIADI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,store_data[11:8]}),
        .DIBDI({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DIPADIP({1'b0,1'b0,1'b0,1'b0}),
        .DIPBDIP({1'b1,1'b1,1'b1,1'b1}),
        .DOADO({NLW_memory_reg_2_DOADO_UNCONNECTED[31:4],load_data[11:8]}),
        .DOBDO(NLW_memory_reg_2_DOBDO_UNCONNECTED[31:0]),
        .DOPADOP(NLW_memory_reg_2_DOPADOP_UNCONNECTED[3:0]),
        .DOPBDOP(NLW_memory_reg_2_DOPBDOP_UNCONNECTED[3:0]),
        .ECCPARITY(NLW_memory_reg_2_ECCPARITY_UNCONNECTED[7:0]),
        .ENARDEN(memory_reg_2_ENARDEN_cooolgate_en_sig_2),
        .ENBWREN(1'b0),
        .INJECTDBITERR(NLW_memory_reg_2_INJECTDBITERR_UNCONNECTED),
        .INJECTSBITERR(NLW_memory_reg_2_INJECTSBITERR_UNCONNECTED),
        .RDADDRECC(NLW_memory_reg_2_RDADDRECC_UNCONNECTED[8:0]),
        .REGCEAREGCE(NLW_memory_reg_2_REGCEAREGCE_UNCONNECTED),
        .REGCEB(NLW_memory_reg_2_REGCEB_UNCONNECTED),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SBITERR(NLW_memory_reg_2_SBITERR_UNCONNECTED),
        .WEA({1'b0,1'b0,1'b0,p_0_in}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
  LUT4 #(
    .INIT(16'hff02))
    memory_reg_2_ENARDEN_cooolgate_en_gate_3
       (.I0(\state[2]_i_1_n_0 ),
        .I1(\state[0]_i_1_n_0 ),
        .I2(INTERNAL_RST_reg),
        .I3(p_0_in),
        .O(memory_reg_2_ENARDEN_cooolgate_en_sig_2));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_2_i_1
       (.I0(result[11]),
        .I1(operand_b1),
        .I2(register_b[11]),
        .O(store_data[11]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_2_i_2
       (.I0(result[10]),
        .I1(operand_b1),
        .I2(register_b[10]),
        .O(store_data[10]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_2_i_3
       (.I0(result[9]),
        .I1(operand_b1),
        .I2(register_b[9]),
        .O(store_data[9]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_2_i_4
       (.I0(result[8]),
        .I1(operand_b1),
        .I2(register_b[8]),
        .O(store_data[8]));
  (* IS_CLOCK_GATED *)
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *)
  (* POWER_OPTED_CE = "ENARDEN=NEW" *)
  (* RTL_RAM_BITS = "131104" *)
  (* RTL_RAM_NAME = "memory" *)
  (* bram_addr_begin = "0" *)
  (* bram_addr_end = "8191" *)
  (* bram_slice_begin = "12" *)
  (* bram_slice_end = "15" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(0))
    memory_reg_3
       (.ADDRARDADDR({1'b1,\write_output[12]_i_1_n_0 ,\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 ,\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 ,\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 ,1'b1,1'b1}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .CASCADEINA(1'b1),
        .CASCADEINB(1'b0),
        .CASCADEOUTA(NLW_memory_reg_3_CASCADEOUTA_UNCONNECTED),
        .CASCADEOUTB(NLW_memory_reg_3_CASCADEOUTB_UNCONNECTED),
        .CLKARDCLK(ETH_CLK_OBUF),
        .CLKBWRCLK(1'b0),
        .DBITERR(NLW_memory_reg_3_DBITERR_UNCONNECTED),
        .DIADI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,store_data[15:12]}),
        .DIBDI({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DIPADIP({1'b0,1'b0,1'b0,1'b0}),
        .DIPBDIP({1'b1,1'b1,1'b1,1'b1}),
        .DOADO({NLW_memory_reg_3_DOADO_UNCONNECTED[31:4],load_data[15:12]}),
        .DOBDO(NLW_memory_reg_3_DOBDO_UNCONNECTED[31:0]),
        .DOPADOP(NLW_memory_reg_3_DOPADOP_UNCONNECTED[3:0]),
        .DOPBDOP(NLW_memory_reg_3_DOPBDOP_UNCONNECTED[3:0]),
        .ECCPARITY(NLW_memory_reg_3_ECCPARITY_UNCONNECTED[7:0]),
        .ENARDEN(memory_reg_3_ENARDEN_cooolgate_en_sig_3),
        .ENBWREN(1'b0),
        .INJECTDBITERR(NLW_memory_reg_3_INJECTDBITERR_UNCONNECTED),
        .INJECTSBITERR(NLW_memory_reg_3_INJECTSBITERR_UNCONNECTED),
        .RDADDRECC(NLW_memory_reg_3_RDADDRECC_UNCONNECTED[8:0]),
        .REGCEAREGCE(NLW_memory_reg_3_REGCEAREGCE_UNCONNECTED),
        .REGCEB(NLW_memory_reg_3_REGCEB_UNCONNECTED),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SBITERR(NLW_memory_reg_3_SBITERR_UNCONNECTED),
        .WEA({1'b0,1'b0,1'b0,p_0_in}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
  LUT4 #(
    .INIT(16'hff02))
    memory_reg_3_ENARDEN_cooolgate_en_gate_5
       (.I0(\state[2]_i_1_n_0 ),
        .I1(\state[0]_i_1_n_0 ),
        .I2(INTERNAL_RST_reg),
        .I3(p_0_in),
        .O(memory_reg_3_ENARDEN_cooolgate_en_sig_3));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_3_i_1
       (.I0(result[15]),
        .I1(operand_b1),
        .I2(register_b[15]),
        .O(store_data[15]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_3_i_2
       (.I0(result[14]),
        .I1(operand_b1),
        .I2(register_b[14]),
        .O(store_data[14]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_3_i_3
       (.I0(result[13]),
        .I1(operand_b1),
        .I2(register_b[13]),
        .O(store_data[13]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_3_i_4
       (.I0(result[12]),
        .I1(operand_b1),
        .I2(register_b[12]),
        .O(store_data[12]));
  (* IS_CLOCK_GATED *)
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *)
  (* POWER_OPTED_CE = "ENARDEN=NEW" *)
  (* RTL_RAM_BITS = "131104" *)
  (* RTL_RAM_NAME = "memory" *)
  (* bram_addr_begin = "0" *)
  (* bram_addr_end = "8191" *)
  (* bram_slice_begin = "16" *)
  (* bram_slice_end = "19" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(0))
    memory_reg_4
       (.ADDRARDADDR({1'b1,\write_output[12]_i_1_n_0 ,\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 ,\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 ,\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 ,1'b1,1'b1}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .CASCADEINA(1'b1),
        .CASCADEINB(1'b0),
        .CASCADEOUTA(NLW_memory_reg_4_CASCADEOUTA_UNCONNECTED),
        .CASCADEOUTB(NLW_memory_reg_4_CASCADEOUTB_UNCONNECTED),
        .CLKARDCLK(ETH_CLK_OBUF),
        .CLKBWRCLK(1'b0),
        .DBITERR(NLW_memory_reg_4_DBITERR_UNCONNECTED),
        .DIADI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,store_data[19:16]}),
        .DIBDI({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DIPADIP({1'b0,1'b0,1'b0,1'b0}),
        .DIPBDIP({1'b1,1'b1,1'b1,1'b1}),
        .DOADO({NLW_memory_reg_4_DOADO_UNCONNECTED[31:4],load_data[19:16]}),
        .DOBDO(NLW_memory_reg_4_DOBDO_UNCONNECTED[31:0]),
        .DOPADOP(NLW_memory_reg_4_DOPADOP_UNCONNECTED[3:0]),
        .DOPBDOP(NLW_memory_reg_4_DOPBDOP_UNCONNECTED[3:0]),
        .ECCPARITY(NLW_memory_reg_4_ECCPARITY_UNCONNECTED[7:0]),
        .ENARDEN(memory_reg_4_ENARDEN_cooolgate_en_sig_4),
        .ENBWREN(1'b0),
        .INJECTDBITERR(NLW_memory_reg_4_INJECTDBITERR_UNCONNECTED),
        .INJECTSBITERR(NLW_memory_reg_4_INJECTSBITERR_UNCONNECTED),
        .RDADDRECC(NLW_memory_reg_4_RDADDRECC_UNCONNECTED[8:0]),
        .REGCEAREGCE(NLW_memory_reg_4_REGCEAREGCE_UNCONNECTED),
        .REGCEB(NLW_memory_reg_4_REGCEB_UNCONNECTED),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SBITERR(NLW_memory_reg_4_SBITERR_UNCONNECTED),
        .WEA({1'b0,1'b0,1'b0,p_0_in}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
  LUT4 #(
    .INIT(16'hff02))
    memory_reg_4_ENARDEN_cooolgate_en_gate_7
       (.I0(\state[2]_i_1_n_0 ),
        .I1(\state[0]_i_1_n_0 ),
        .I2(INTERNAL_RST_reg),
        .I3(p_0_in),
        .O(memory_reg_4_ENARDEN_cooolgate_en_sig_4));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_4_i_1
       (.I0(result[19]),
        .I1(operand_b1),
        .I2(register_b[19]),
        .O(store_data[19]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_4_i_2
       (.I0(result[18]),
        .I1(operand_b1),
        .I2(register_b[18]),
        .O(store_data[18]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_4_i_3
       (.I0(result[17]),
        .I1(operand_b1),
        .I2(register_b[17]),
        .O(store_data[17]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_4_i_4
       (.I0(result[16]),
        .I1(operand_b1),
        .I2(register_b[16]),
        .O(store_data[16]));
  (* IS_CLOCK_GATED *)
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *)
  (* POWER_OPTED_CE = "ENARDEN=NEW" *)
  (* RTL_RAM_BITS = "131104" *)
  (* RTL_RAM_NAME = "memory" *)
  (* bram_addr_begin = "0" *)
  (* bram_addr_end = "8191" *)
  (* bram_slice_begin = "20" *)
  (* bram_slice_end = "23" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(0))
    memory_reg_5
       (.ADDRARDADDR({1'b1,\write_output[12]_i_1_n_0 ,\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 ,\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 ,\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 ,1'b1,1'b1}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .CASCADEINA(1'b1),
        .CASCADEINB(1'b0),
        .CASCADEOUTA(NLW_memory_reg_5_CASCADEOUTA_UNCONNECTED),
        .CASCADEOUTB(NLW_memory_reg_5_CASCADEOUTB_UNCONNECTED),
        .CLKARDCLK(ETH_CLK_OBUF),
        .CLKBWRCLK(1'b0),
        .DBITERR(NLW_memory_reg_5_DBITERR_UNCONNECTED),
        .DIADI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,store_data[23:20]}),
        .DIBDI({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DIPADIP({1'b0,1'b0,1'b0,1'b0}),
        .DIPBDIP({1'b1,1'b1,1'b1,1'b1}),
        .DOADO({NLW_memory_reg_5_DOADO_UNCONNECTED[31:4],load_data[23:20]}),
        .DOBDO(NLW_memory_reg_5_DOBDO_UNCONNECTED[31:0]),
        .DOPADOP(NLW_memory_reg_5_DOPADOP_UNCONNECTED[3:0]),
        .DOPBDOP(NLW_memory_reg_5_DOPBDOP_UNCONNECTED[3:0]),
        .ECCPARITY(NLW_memory_reg_5_ECCPARITY_UNCONNECTED[7:0]),
        .ENARDEN(memory_reg_5_ENARDEN_cooolgate_en_sig_5),
        .ENBWREN(1'b0),
        .INJECTDBITERR(NLW_memory_reg_5_INJECTDBITERR_UNCONNECTED),
        .INJECTSBITERR(NLW_memory_reg_5_INJECTSBITERR_UNCONNECTED),
        .RDADDRECC(NLW_memory_reg_5_RDADDRECC_UNCONNECTED[8:0]),
        .REGCEAREGCE(NLW_memory_reg_5_REGCEAREGCE_UNCONNECTED),
        .REGCEB(NLW_memory_reg_5_REGCEB_UNCONNECTED),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SBITERR(NLW_memory_reg_5_SBITERR_UNCONNECTED),
        .WEA({1'b0,1'b0,1'b0,p_0_in}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
  LUT4 #(
    .INIT(16'hff02))
    memory_reg_5_ENARDEN_cooolgate_en_gate_9
       (.I0(\state[2]_i_1_n_0 ),
        .I1(\state[0]_i_1_n_0 ),
        .I2(INTERNAL_RST_reg),
        .I3(p_0_in),
        .O(memory_reg_5_ENARDEN_cooolgate_en_sig_5));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_5_i_1
       (.I0(result[23]),
        .I1(operand_b1),
        .I2(register_b[23]),
        .O(store_data[23]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_5_i_2
       (.I0(result[22]),
        .I1(operand_b1),
        .I2(register_b[22]),
        .O(store_data[22]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_5_i_3
       (.I0(result[21]),
        .I1(operand_b1),
        .I2(register_b[21]),
        .O(store_data[21]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_5_i_4
       (.I0(result[20]),
        .I1(operand_b1),
        .I2(register_b[20]),
        .O(store_data[20]));
  (* IS_CLOCK_GATED *)
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *)
  (* POWER_OPTED_CE = "ENARDEN=NEW" *)
  (* RTL_RAM_BITS = "131104" *)
  (* RTL_RAM_NAME = "memory" *)
  (* bram_addr_begin = "0" *)
  (* bram_addr_end = "8191" *)
  (* bram_slice_begin = "24" *)
  (* bram_slice_end = "27" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(0))
    memory_reg_6
       (.ADDRARDADDR({1'b1,\write_output[12]_i_1_n_0 ,\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 ,\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 ,\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 ,1'b1,1'b1}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .CASCADEINA(1'b1),
        .CASCADEINB(1'b0),
        .CASCADEOUTA(NLW_memory_reg_6_CASCADEOUTA_UNCONNECTED),
        .CASCADEOUTB(NLW_memory_reg_6_CASCADEOUTB_UNCONNECTED),
        .CLKARDCLK(ETH_CLK_OBUF),
        .CLKBWRCLK(1'b0),
        .DBITERR(NLW_memory_reg_6_DBITERR_UNCONNECTED),
        .DIADI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,store_data[27:24]}),
        .DIBDI({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DIPADIP({1'b0,1'b0,1'b0,1'b0}),
        .DIPBDIP({1'b1,1'b1,1'b1,1'b1}),
        .DOADO({NLW_memory_reg_6_DOADO_UNCONNECTED[31:4],load_data[27:24]}),
        .DOBDO(NLW_memory_reg_6_DOBDO_UNCONNECTED[31:0]),
        .DOPADOP(NLW_memory_reg_6_DOPADOP_UNCONNECTED[3:0]),
        .DOPBDOP(NLW_memory_reg_6_DOPBDOP_UNCONNECTED[3:0]),
        .ECCPARITY(NLW_memory_reg_6_ECCPARITY_UNCONNECTED[7:0]),
        .ENARDEN(memory_reg_6_ENARDEN_cooolgate_en_sig_6),
        .ENBWREN(1'b0),
        .INJECTDBITERR(NLW_memory_reg_6_INJECTDBITERR_UNCONNECTED),
        .INJECTSBITERR(NLW_memory_reg_6_INJECTSBITERR_UNCONNECTED),
        .RDADDRECC(NLW_memory_reg_6_RDADDRECC_UNCONNECTED[8:0]),
        .REGCEAREGCE(NLW_memory_reg_6_REGCEAREGCE_UNCONNECTED),
        .REGCEB(NLW_memory_reg_6_REGCEB_UNCONNECTED),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SBITERR(NLW_memory_reg_6_SBITERR_UNCONNECTED),
        .WEA({1'b0,1'b0,1'b0,p_0_in}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
  LUT4 #(
    .INIT(16'hff02))
    memory_reg_6_ENARDEN_cooolgate_en_gate_11
       (.I0(\state[2]_i_1_n_0 ),
        .I1(\state[0]_i_1_n_0 ),
        .I2(INTERNAL_RST_reg),
        .I3(p_0_in),
        .O(memory_reg_6_ENARDEN_cooolgate_en_sig_6));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_6_i_1
       (.I0(result[27]),
        .I1(operand_b1),
        .I2(register_b[27]),
        .O(store_data[27]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_6_i_2
       (.I0(result[26]),
        .I1(operand_b1),
        .I2(register_b[26]),
        .O(store_data[26]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_6_i_3
       (.I0(result[25]),
        .I1(operand_b1),
        .I2(register_b[25]),
        .O(store_data[25]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_6_i_4
       (.I0(result[24]),
        .I1(operand_b1),
        .I2(register_b[24]),
        .O(store_data[24]));
  (* IS_CLOCK_GATED *)
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *)
  (* POWER_OPTED_CE = "ENARDEN=NEW" *)
  (* RTL_RAM_BITS = "131104" *)
  (* RTL_RAM_NAME = "memory" *)
  (* bram_addr_begin = "0" *)
  (* bram_addr_end = "8191" *)
  (* bram_slice_begin = "28" *)
  (* bram_slice_end = "31" *)
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(4),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(4),
    .WRITE_WIDTH_B(0))
    memory_reg_7
       (.ADDRARDADDR({1'b1,\write_output[12]_i_1_n_0 ,\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 ,\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 ,\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 ,1'b1,1'b1}),
        .ADDRBWRADDR({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .CASCADEINA(1'b1),
        .CASCADEINB(1'b0),
        .CASCADEOUTA(NLW_memory_reg_7_CASCADEOUTA_UNCONNECTED),
        .CASCADEOUTB(NLW_memory_reg_7_CASCADEOUTB_UNCONNECTED),
        .CLKARDCLK(ETH_CLK_OBUF),
        .CLKBWRCLK(1'b0),
        .DBITERR(NLW_memory_reg_7_DBITERR_UNCONNECTED),
        .DIADI({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,store_data[31:28]}),
        .DIBDI({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),
        .DIPADIP({1'b0,1'b0,1'b0,1'b0}),
        .DIPBDIP({1'b1,1'b1,1'b1,1'b1}),
        .DOADO({NLW_memory_reg_7_DOADO_UNCONNECTED[31:4],load_data[31:28]}),
        .DOBDO(NLW_memory_reg_7_DOBDO_UNCONNECTED[31:0]),
        .DOPADOP(NLW_memory_reg_7_DOPADOP_UNCONNECTED[3:0]),
        .DOPBDOP(NLW_memory_reg_7_DOPBDOP_UNCONNECTED[3:0]),
        .ECCPARITY(NLW_memory_reg_7_ECCPARITY_UNCONNECTED[7:0]),
        .ENARDEN(memory_reg_7_ENARDEN_cooolgate_en_sig_7),
        .ENBWREN(1'b0),
        .INJECTDBITERR(NLW_memory_reg_7_INJECTDBITERR_UNCONNECTED),
        .INJECTSBITERR(NLW_memory_reg_7_INJECTSBITERR_UNCONNECTED),
        .RDADDRECC(NLW_memory_reg_7_RDADDRECC_UNCONNECTED[8:0]),
        .REGCEAREGCE(NLW_memory_reg_7_REGCEAREGCE_UNCONNECTED),
        .REGCEB(NLW_memory_reg_7_REGCEB_UNCONNECTED),
        .RSTRAMARSTRAM(1'b0),
        .RSTRAMB(1'b0),
        .RSTREGARSTREG(1'b0),
        .RSTREGB(1'b0),
        .SBITERR(NLW_memory_reg_7_SBITERR_UNCONNECTED),
        .WEA({1'b0,1'b0,1'b0,p_0_in}),
        .WEBWE({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
  LUT4 #(
    .INIT(16'hff02))
    memory_reg_7_ENARDEN_cooolgate_en_gate_13
       (.I0(\state[2]_i_1_n_0 ),
        .I1(\state[0]_i_1_n_0 ),
        .I2(INTERNAL_RST_reg),
        .I3(p_0_in),
        .O(memory_reg_7_ENARDEN_cooolgate_en_sig_7));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_7_i_1
       (.I0(result[31]),
        .I1(operand_b1),
        .I2(register_b[31]),
        .O(store_data[31]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_7_i_2
       (.I0(result[30]),
        .I1(operand_b1),
        .I2(register_b[30]),
        .O(store_data[30]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_7_i_3
       (.I0(result[29]),
        .I1(operand_b1),
        .I2(register_b[29]),
        .O(store_data[29]));
  LUT3 #(
    .INIT(8'hB8))
    memory_reg_7_i_4
       (.I0(result[28]),
        .I1(operand_b1),
        .I2(register_b[28]),
        .O(store_data[28]));
  LUT2 #(
    .INIT(4'h2))
    \opcode_2[3]_i_1
       (.I0(\state_reg_n_0_[1] ),
        .I1(\state_reg_n_0_[2] ),
        .O(opcode_20));
  FDRE \opcode_2_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(opcode[0]),
        .Q(opcode_2[0]),
        .R(1'b0));
  FDRE \opcode_2_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(opcode[1]),
        .Q(opcode_2[1]),
        .R(1'b0));
  FDRE \opcode_2_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(opcode[2]),
        .Q(opcode_2[2]),
        .R(1'b0));
  FDRE \opcode_2_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(opcode[3]),
        .Q(opcode_2[3]),
        .R(1'b0));
  LUT5 #(
    .INIT(32'hFFEAEAEA))
    \program_counter[10]_i_1
       (.I0(\program_counter[15]_i_2_n_0 ),
        .I1(\program_counter_rep[9]_i_4_n_0 ),
        .I2(data1[10]),
        .I3(\write_output[10]_i_1_n_0 ),
        .I4(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter[10]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA))
    \program_counter[11]_i_1
       (.I0(\program_counter[15]_i_2_n_0 ),
        .I1(\program_counter_rep[9]_i_4_n_0 ),
        .I2(data1[11]),
        .I3(\write_output[11]_i_1_n_0 ),
        .I4(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA))
    \program_counter[12]_i_1
       (.I0(\program_counter[15]_i_2_n_0 ),
        .I1(\program_counter_rep[9]_i_6_n_0 ),
        .I2(\write_output[12]_i_1_n_0 ),
        .I3(data1[12]),
        .I4(\program_counter_rep[9]_i_4_n_0 ),
        .O(\program_counter[12]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA))
    \program_counter[13]_i_1
       (.I0(\program_counter[15]_i_2_n_0 ),
        .I1(\program_counter_rep[9]_i_6_n_0 ),
        .I2(\write_output[13]_i_1_n_0 ),
        .I3(data1[13]),
        .I4(\program_counter_rep[9]_i_4_n_0 ),
        .O(\program_counter[13]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA))
    \program_counter[14]_i_1
       (.I0(\program_counter[15]_i_2_n_0 ),
        .I1(\program_counter_rep[9]_i_6_n_0 ),
        .I2(\write_output[14]_i_1_n_0 ),
        .I3(data1[14]),
        .I4(\program_counter_rep[9]_i_4_n_0 ),
        .O(\program_counter[14]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA))
    \program_counter[15]_i_1
       (.I0(\program_counter[15]_i_2_n_0 ),
        .I1(\program_counter_rep[9]_i_6_n_0 ),
        .I2(\write_output[15]_i_1_n_0 ),
        .I3(data1[15]),
        .I4(\program_counter_rep[9]_i_4_n_0 ),
        .O(\program_counter[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE))
    \program_counter[15]_i_11
       (.I0(\write_output[21]_i_1_n_0 ),
        .I1(\program_counter[15]_i_13_n_0 ),
        .I2(\program_counter[15]_i_14_n_0 ),
        .I3(\write_output[27]_i_1_n_0 ),
        .I4(\program_counter[15]_i_15_n_0 ),
        .I5(\write_output[24]_i_1_n_0 ),
        .O(\program_counter[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE))
    \program_counter[15]_i_12
       (.I0(\write_output[12]_i_1_n_0 ),
        .I1(\program_counter[15]_i_16_n_0 ),
        .I2(\program_counter[15]_i_17_n_0 ),
        .I3(\write_output[3]_i_1_n_0 ),
        .I4(\program_counter[15]_i_18_n_0 ),
        .I5(\write_output[0]_i_1_n_0 ),
        .O(\program_counter[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAFAFACCFAFAFA))
    \program_counter[15]_i_13
       (.I0(register_a[22]),
        .I1(result[22]),
        .I2(register_a[23]),
        .I3(\program_counter_rep[9]_i_22_n_0 ),
        .I4(\write_output[31]_i_4_n_0 ),
        .I5(result[23]),
        .O(\program_counter[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAFAFACCFAFAFA))
    \program_counter[15]_i_14
       (.I0(register_a[28]),
        .I1(result[28]),
        .I2(register_a[29]),
        .I3(\program_counter_rep[9]_i_22_n_0 ),
        .I4(\write_output[31]_i_4_n_0 ),
        .I5(result[29]),
        .O(\program_counter[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAFAFACCFAFAFA))
    \program_counter[15]_i_15
       (.I0(register_a[25]),
        .I1(result[25]),
        .I2(register_a[26]),
        .I3(\program_counter_rep[9]_i_22_n_0 ),
        .I4(\write_output[31]_i_4_n_0 ),
        .I5(result[26]),
        .O(\program_counter[15]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAFAFACCFAFAFA))
    \program_counter[15]_i_16
       (.I0(register_a[13]),
        .I1(result[13]),
        .I2(register_a[14]),
        .I3(\program_counter_rep[9]_i_22_n_0 ),
        .I4(\write_output[31]_i_4_n_0 ),
        .I5(result[14]),
        .O(\program_counter[15]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAFAFACCFAFAFA))
    \program_counter[15]_i_17
       (.I0(register_a[4]),
        .I1(result[4]),
        .I2(register_a[5]),
        .I3(\program_counter_rep[9]_i_22_n_0 ),
        .I4(\write_output[31]_i_4_n_0 ),
        .I5(result[5]),
        .O(\program_counter[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAFAFACCFAFAFA))
    \program_counter[15]_i_18
       (.I0(register_a[1]),
        .I1(result[1]),
        .I2(register_a[2]),
        .I3(\program_counter_rep[9]_i_22_n_0 ),
        .I4(\write_output[31]_i_4_n_0 ),
        .I5(result[2]),
        .O(\program_counter[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFF8F8F8F0F0F0F0))
    \program_counter[15]_i_2
       (.I0(\program_counter_rep[9]_i_7_n_0 ),
        .I1(\program_counter[15]_i_4_n_0 ),
        .I2(\program_counter[15]_i_5_n_0 ),
        .I3(\program_counter[15]_i_6_n_0 ),
        .I4(\program_counter[15]_i_7_n_0 ),
        .I5(literal_2[15]),
        .O(\program_counter[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000))
    \program_counter[15]_i_4
       (.I0(opcode_2[3]),
        .I1(\state_reg_n_0_[1] ),
        .I2(opcode_2[1]),
        .I3(opcode_2[0]),
        .I4(opcode_2[2]),
        .I5(\state_reg_n_0_[0] ),
        .O(\program_counter[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h80000000))
    \program_counter[15]_i_5
       (.I0(literal_2[15]),
        .I1(memory_reg_0_i_2_n_0),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(\state_reg_n_0_[1] ),
        .O(\program_counter[15]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0800))
    \program_counter[15]_i_6
       (.I0(\state_reg_n_0_[1] ),
        .I1(opcode_2[3]),
        .I2(opcode_2[2]),
        .I3(\state_reg_n_0_[0] ),
        .O(\program_counter[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0001))
    \program_counter[15]_i_7
       (.I0(\program_counter[15]_i_11_n_0 ),
        .I1(\program_counter_rep[9]_i_16_n_0 ),
        .I2(\program_counter_rep[9]_i_17_n_0 ),
        .I3(\program_counter[15]_i_12_n_0 ),
        .I4(opcode_2[0]),
        .I5(opcode_2[1]),
        .O(\program_counter[15]_i_7_n_0 ));
  FDRE \program_counter_1_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[0] ),
        .Q(program_counter_1[0]),
        .R(1'b0));
  FDRE \program_counter_1_reg[10]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[10] ),
        .Q(program_counter_1[10]),
        .R(1'b0));
  FDRE \program_counter_1_reg[11]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[11] ),
        .Q(program_counter_1[11]),
        .R(1'b0));
  FDRE \program_counter_1_reg[12]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[12] ),
        .Q(program_counter_1[12]),
        .R(1'b0));
  FDRE \program_counter_1_reg[13]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[13] ),
        .Q(program_counter_1[13]),
        .R(1'b0));
  FDRE \program_counter_1_reg[14]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[14] ),
        .Q(program_counter_1[14]),
        .R(1'b0));
  FDRE \program_counter_1_reg[15]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[15] ),
        .Q(program_counter_1[15]),
        .R(1'b0));
  FDRE \program_counter_1_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[1] ),
        .Q(program_counter_1[1]),
        .R(1'b0));
  FDRE \program_counter_1_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[2] ),
        .Q(program_counter_1[2]),
        .R(1'b0));
  FDRE \program_counter_1_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[3] ),
        .Q(program_counter_1[3]),
        .R(1'b0));
  FDRE \program_counter_1_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[4] ),
        .Q(program_counter_1[4]),
        .R(1'b0));
  FDRE \program_counter_1_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[5] ),
        .Q(program_counter_1[5]),
        .R(1'b0));
  FDRE \program_counter_1_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[6] ),
        .Q(program_counter_1[6]),
        .R(1'b0));
  FDRE \program_counter_1_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[7] ),
        .Q(program_counter_1[7]),
        .R(1'b0));
  FDRE \program_counter_1_reg[8]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[8] ),
        .Q(program_counter_1[8]),
        .R(1'b0));
  FDRE \program_counter_1_reg[9]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_reg_n_0_[9] ),
        .Q(program_counter_1[9]),
        .R(1'b0));
  FDRE \program_counter_2_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[0]),
        .Q(program_counter_2[0]),
        .R(1'b0));
  FDRE \program_counter_2_reg[10]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[10]),
        .Q(program_counter_2[10]),
        .R(1'b0));
  FDRE \program_counter_2_reg[11]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[11]),
        .Q(program_counter_2[11]),
        .R(1'b0));
  FDRE \program_counter_2_reg[12]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[12]),
        .Q(program_counter_2[12]),
        .R(1'b0));
  FDRE \program_counter_2_reg[13]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[13]),
        .Q(program_counter_2[13]),
        .R(1'b0));
  FDRE \program_counter_2_reg[14]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[14]),
        .Q(program_counter_2[14]),
        .R(1'b0));
  FDRE \program_counter_2_reg[15]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[15]),
        .Q(program_counter_2[15]),
        .R(1'b0));
  FDRE \program_counter_2_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[1]),
        .Q(program_counter_2[1]),
        .R(1'b0));
  FDRE \program_counter_2_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[2]),
        .Q(program_counter_2[2]),
        .R(1'b0));
  FDRE \program_counter_2_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[3]),
        .Q(program_counter_2[3]),
        .R(1'b0));
  FDRE \program_counter_2_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[4]),
        .Q(program_counter_2[4]),
        .R(1'b0));
  FDRE \program_counter_2_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[5]),
        .Q(program_counter_2[5]),
        .R(1'b0));
  FDRE \program_counter_2_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[6]),
        .Q(program_counter_2[6]),
        .R(1'b0));
  FDRE \program_counter_2_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[7]),
        .Q(program_counter_2[7]),
        .R(1'b0));
  FDRE \program_counter_2_reg[8]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[8]),
        .Q(program_counter_2[8]),
        .R(1'b0));
  FDRE \program_counter_2_reg[9]
       (.C(ETH_CLK_OBUF),
        .CE(opcode_20),
        .D(program_counter_1[9]),
        .Q(program_counter_2[9]),
        .R(1'b0));
  FDRE \program_counter_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[0]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[0] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[10]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter[10]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[10] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[11]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter[11]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[11] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[12]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter[12]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[12] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[13]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter[13]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[13] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[14]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter[14]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[14] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[15]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter[15]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[15] ),
        .R(INTERNAL_RST_reg));
  CARRY4 \program_counter_reg[15]_i_3
       (.CI(\program_counter_reg_rep[9]_i_5_n_0 ),
        .CO(\NLW_program_counter_reg[15]_i_3_CO_UNCONNECTED [3:0]),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_program_counter_reg[15]_i_3_O_UNCONNECTED [3],data1[15:13]}),
        .S({1'b0,\program_counter_reg_n_0_[15] ,\program_counter_reg_n_0_[14] ,\program_counter_reg_n_0_[13] }));
  FDRE \program_counter_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[1]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[1] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[2]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[2] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[3]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[3] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[4]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[4] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[5]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[5] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[6]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[6] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[7]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[7] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[8]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[8]_i_1_n_0 ),
        .Q(\program_counter_reg_n_0_[8] ),
        .R(INTERNAL_RST_reg));
  FDRE \program_counter_reg[9]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[9]_i_2_n_0 ),
        .Q(\program_counter_reg_n_0_[9] ),
        .R(INTERNAL_RST_reg));
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[0]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[0]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[0] ),
        .R(INTERNAL_RST_reg));
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[1]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[1]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[1] ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[2]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[2]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[2]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[2] ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[2]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[2]_rep
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[2]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[2]_rep_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[2]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[2]_rep__0
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[2]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[2]_rep__0_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[3]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[3]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[3]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[3] ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[3]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[3]_rep
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[3]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[3]_rep_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[3]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[3]_rep__0
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[3]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[3]_rep__0_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[3]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[3]_rep__1
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[3]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[3]_rep__1_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[4]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[4]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[4]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[4] ),
        .R(INTERNAL_RST_reg));
  CARRY4 \program_counter_reg_rep[4]_i_2
       (.CI(1'b0),
        .CO({\program_counter_reg_rep[4]_i_2_n_0 ,\NLW_program_counter_reg_rep[4]_i_2_CO_UNCONNECTED [2:0]}),
        .CYINIT(\program_counter_reg_n_0_[0] ),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(data1[4:1]),
        .S({\program_counter_reg_n_0_[4] ,\program_counter_reg_n_0_[3] ,\program_counter_reg_n_0_[2] ,\program_counter_reg_n_0_[1] }));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[4]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[4]_rep
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[4]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[4]_rep_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[4]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[4]_rep__0
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[4]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[4]_rep__0_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[4]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[4]_rep__1
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[4]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[4]_rep__1_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[4]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[4]_rep__2
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[4]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[4]_rep__2_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[5]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[5]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[5]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[5] ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[5]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[5]_rep
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[5]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[5]_rep_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[5]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[5]_rep__0
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[5]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[5]_rep__0_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[5]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[5]_rep__1
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[5]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[5]_rep__1_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[5]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[5]_rep__2
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[5]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[5]_rep__2_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[6]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[6]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[6]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[6] ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[6]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[6]_rep
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[6]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[6]_rep_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[6]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[6]_rep__0
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[6]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[6]_rep__0_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[6]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[6]_rep__1
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[6]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[6]_rep__1_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[6]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[6]_rep__2
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[6]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[6]_rep__2_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[7]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[7]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[7]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[7] ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[7]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[7]_rep
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[7]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[7]_rep_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[7]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[7]_rep__0
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[7]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[7]_rep__0_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[7]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[7]_rep__1
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[7]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[7]_rep__1_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[8]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[8]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[8]_i_1_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[8] ),
        .R(INTERNAL_RST_reg));
  CARRY4 \program_counter_reg_rep[8]_i_2
       (.CI(\program_counter_reg_rep[4]_i_2_n_0 ),
        .CO({\program_counter_reg_rep[8]_i_2_n_0 ,\NLW_program_counter_reg_rep[8]_i_2_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(data1[8:5]),
        .S({\program_counter_reg_n_0_[8] ,\program_counter_reg_n_0_[7] ,\program_counter_reg_n_0_[6] ,\program_counter_reg_n_0_[5] }));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[8]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[8]_rep
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[8]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[8]_rep_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[8]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[8]_rep__0
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[8]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[8]_rep__0_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[8]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[8]_rep__1
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[8]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[8]_rep__1_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[8]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[8]_rep__2
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[8]_i_1_n_0 ),
        .Q(\program_counter_reg_rep[8]_rep__2_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[9]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[9]
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[9]_i_2_n_0 ),
        .Q(\program_counter_reg_rep_n_0_[9] ),
        .R(INTERNAL_RST_reg));
  CARRY4 \program_counter_reg_rep[9]_i_5
       (.CI(\program_counter_reg_rep[8]_i_2_n_0 ),
        .CO({\program_counter_reg_rep[9]_i_5_n_0 ,\NLW_program_counter_reg_rep[9]_i_5_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(data1[12:9]),
        .S({\program_counter_reg_n_0_[12] ,\program_counter_reg_n_0_[11] ,\program_counter_reg_n_0_[10] ,\program_counter_reg_n_0_[9] }));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[9]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[9]_rep
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[9]_i_2_n_0 ),
        .Q(\program_counter_reg_rep[9]_rep_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[9]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[9]_rep__0
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[9]_i_2_n_0 ),
        .Q(\program_counter_reg_rep[9]_rep__0_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[9]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[9]_rep__1
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[9]_i_2_n_0 ),
        .Q(\program_counter_reg_rep[9]_rep__1_n_0 ),
        .R(INTERNAL_RST_reg));
  (* ORIG_CELL_NAME = "program_counter_reg_rep[9]" *)
  (* equivalent_register_removal = "no" *)
  FDRE \program_counter_reg_rep[9]_rep__2
       (.C(ETH_CLK_OBUF),
        .CE(instruction0),
        .D(\program_counter_rep[9]_i_2_n_0 ),
        .Q(\program_counter_reg_rep[9]_rep__2_n_0 ),
        .R(INTERNAL_RST_reg));
  LUT6 #(
    .INIT(64'hFFFFF222F222F222))
    \program_counter_rep[0]_i_1
       (.I0(\program_counter_rep[9]_i_4_n_0 ),
        .I1(\program_counter_reg_n_0_[0] ),
        .I2(\program_counter_rep[9]_i_6_n_0 ),
        .I3(\write_output[0]_i_1_n_0 ),
        .I4(address_b_2[0]),
        .I5(\program_counter_rep[9]_i_3_n_0 ),
        .O(\program_counter_rep[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[1]_i_1
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(address_b_2[1]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[1]),
        .I4(\write_output[1]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[2]_i_1
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(address_b_2[2]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[2]),
        .I4(\write_output[2]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[3]_i_1
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(address_b_2[3]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[3]),
        .I4(\write_output[3]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[4]_i_1
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(literal_2[4]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[4]),
        .I4(\write_output[4]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[5]_i_1
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(literal_2[5]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[5]),
        .I4(\write_output[5]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[6]_i_1
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(literal_2[6]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[6]),
        .I4(\write_output[6]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[7]_i_1
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(literal_2[7]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[7]),
        .I4(\write_output[7]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[8]_i_1
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(literal_2[8]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[8]),
        .I4(\write_output[8]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h0E))
    \program_counter_rep[9]_i_1
       (.I0(\state_reg_n_0_[1] ),
        .I1(\state_reg_n_0_[0] ),
        .I2(\state_reg_n_0_[2] ),
        .O(instruction0));
  LUT6 #(
    .INIT(64'hFFFFFFFCFAFAFFFC))
    \program_counter_rep[9]_i_14
       (.I0(result[23]),
        .I1(register_a[23]),
        .I2(\write_output[22]_i_1_n_0 ),
        .I3(register_a[21]),
        .I4(operand_a1),
        .I5(result[21]),
        .O(\program_counter_rep[9]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE))
    \program_counter_rep[9]_i_15
       (.I0(\write_output[24]_i_1_n_0 ),
        .I1(\write_output[25]_i_1_n_0 ),
        .I2(\write_output[26]_i_1_n_0 ),
        .I3(\write_output[27]_i_1_n_0 ),
        .I4(\write_output[28]_i_1_n_0 ),
        .I5(\write_output[29]_i_1_n_0 ),
        .O(\program_counter_rep[9]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE))
    \program_counter_rep[9]_i_16
       (.I0(\write_output[15]_i_1_n_0 ),
        .I1(\write_output[16]_i_1_n_0 ),
        .I2(\write_output[17]_i_1_n_0 ),
        .I3(\write_output[18]_i_1_n_0 ),
        .I4(\write_output[19]_i_1_n_0 ),
        .I5(\write_output[20]_i_1_n_0 ),
        .O(\program_counter_rep[9]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE))
    \program_counter_rep[9]_i_17
       (.I0(\write_output[6]_i_1_n_0 ),
        .I1(\write_output[7]_i_1_n_0 ),
        .I2(\write_output[8]_i_1_n_0 ),
        .I3(\program_counter_rep[9]_i_20_n_0 ),
        .I4(\program_counter_rep[9]_i_21_n_0 ),
        .I5(\write_output[9]_i_1_n_0 ),
        .O(\program_counter_rep[9]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBBFCB8))
    \program_counter_rep[9]_i_18
       (.I0(result[14]),
        .I1(operand_a1),
        .I2(register_a[14]),
        .I3(result[13]),
        .I4(register_a[13]),
        .I5(\write_output[12]_i_1_n_0 ),
        .O(\program_counter_rep[9]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE))
    \program_counter_rep[9]_i_19
       (.I0(\write_output[0]_i_1_n_0 ),
        .I1(\write_output[1]_i_1_n_0 ),
        .I2(\write_output[2]_i_1_n_0 ),
        .I3(\write_output[3]_i_1_n_0 ),
        .I4(\write_output[4]_i_1_n_0 ),
        .I5(\write_output[5]_i_1_n_0 ),
        .O(\program_counter_rep[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \program_counter_rep[9]_i_2
       (.I0(\program_counter_rep[9]_i_3_n_0 ),
        .I1(literal_2[9]),
        .I2(\program_counter_rep[9]_i_4_n_0 ),
        .I3(data1[9]),
        .I4(\write_output[9]_i_1_n_0 ),
        .I5(\program_counter_rep[9]_i_6_n_0 ),
        .O(\program_counter_rep[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAFAFACCFAFAFA))
    \program_counter_rep[9]_i_20
       (.I0(register_a[30]),
        .I1(result[30]),
        .I2(register_a[31]),
        .I3(\program_counter_rep[9]_i_22_n_0 ),
        .I4(\write_output[31]_i_4_n_0 ),
        .I5(result[31]),
        .O(\program_counter_rep[9]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAFAFACCFAFAFA))
    \program_counter_rep[9]_i_21
       (.I0(register_a[10]),
        .I1(result[10]),
        .I2(register_a[11]),
        .I3(\program_counter_rep[9]_i_22_n_0 ),
        .I4(\write_output[31]_i_4_n_0 ),
        .I5(result[11]),
        .O(\program_counter_rep[9]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h90))
    \program_counter_rep[9]_i_22
       (.I0(address_z_3[3]),
        .I1(address_a_2[3]),
        .I2(write_enable),
        .O(\program_counter_rep[9]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h08C40000C0000000))
    \program_counter_rep[9]_i_3
       (.I0(\program_counter_rep[9]_i_7_n_0 ),
        .I1(\program_counter_rep[9]_i_8_n_0 ),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(\state_reg_n_0_[1] ),
        .I5(opcode_2[3]),
        .O(\program_counter_rep[9]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hABBA))
    \program_counter_rep[9]_i_4
       (.I0(\program_counter_rep[9]_i_9_n_0 ),
        .I1(opcode_2[0]),
        .I2(opcode_2[1]),
        .I3(\program_counter_rep[9]_i_7_n_0 ),
        .O(\program_counter_rep[9]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000))
    \program_counter_rep[9]_i_6
       (.I0(opcode_2[2]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[3]),
        .I3(\state_reg_n_0_[1] ),
        .I4(opcode_2[0]),
        .I5(opcode_2[1]),
        .O(\program_counter_rep[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE))
    \program_counter_rep[9]_i_7
       (.I0(\program_counter_rep[9]_i_14_n_0 ),
        .I1(\program_counter_rep[9]_i_15_n_0 ),
        .I2(\program_counter_rep[9]_i_16_n_0 ),
        .I3(\program_counter_rep[9]_i_17_n_0 ),
        .I4(\program_counter_rep[9]_i_18_n_0 ),
        .I5(\program_counter_rep[9]_i_19_n_0 ),
        .O(\program_counter_rep[9]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2))
    \program_counter_rep[9]_i_8
       (.I0(\state_reg_n_0_[0] ),
        .I1(opcode_2[2]),
        .O(\program_counter_rep[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FFFDF7F7F7F))
    \program_counter_rep[9]_i_9
       (.I0(\state_reg_n_0_[0] ),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[1] ),
        .I3(opcode_2[0]),
        .I4(opcode_2[1]),
        .I5(opcode_2[2]),
        .O(\program_counter_rep[9]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080))
    \read_input[31]_i_1
       (.I0(opcode_2[2]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[1]),
        .I3(opcode_2[0]),
        .I4(opcode_2[3]),
        .I5(\read_input[31]_i_2_n_0 ),
        .O(\read_input[31]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB))
    \read_input[31]_i_2
       (.I0(\state_reg_n_0_[2] ),
        .I1(\state_reg_n_0_[1] ),
        .O(\read_input[31]_i_2_n_0 ));
  FDRE \read_input_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[0]_i_1_n_0 ),
        .Q(read_input[0]),
        .R(1'b0));
  FDRE \read_input_reg[10]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[10]_i_1_n_0 ),
        .Q(read_input[10]),
        .R(1'b0));
  FDRE \read_input_reg[11]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[11]_i_1_n_0 ),
        .Q(read_input[11]),
        .R(1'b0));
  FDRE \read_input_reg[12]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[12]_i_1_n_0 ),
        .Q(read_input[12]),
        .R(1'b0));
  FDRE \read_input_reg[13]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[13]_i_1_n_0 ),
        .Q(read_input[13]),
        .R(1'b0));
  FDRE \read_input_reg[14]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[14]_i_1_n_0 ),
        .Q(read_input[14]),
        .R(1'b0));
  FDRE \read_input_reg[15]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[15]_i_1_n_0 ),
        .Q(read_input[15]),
        .R(1'b0));
  FDRE \read_input_reg[16]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[16]_i_1_n_0 ),
        .Q(read_input[16]),
        .R(1'b0));
  FDRE \read_input_reg[17]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[17]_i_1_n_0 ),
        .Q(read_input[17]),
        .R(1'b0));
  FDRE \read_input_reg[18]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[18]_i_1_n_0 ),
        .Q(read_input[18]),
        .R(1'b0));
  FDRE \read_input_reg[19]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[19]_i_1_n_0 ),
        .Q(read_input[19]),
        .R(1'b0));
  FDRE \read_input_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[1]_i_1_n_0 ),
        .Q(read_input[1]),
        .R(1'b0));
  FDRE \read_input_reg[20]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[20]_i_1_n_0 ),
        .Q(read_input[20]),
        .R(1'b0));
  FDRE \read_input_reg[21]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[21]_i_1_n_0 ),
        .Q(read_input[21]),
        .R(1'b0));
  FDRE \read_input_reg[22]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[22]_i_1_n_0 ),
        .Q(read_input[22]),
        .R(1'b0));
  FDRE \read_input_reg[23]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[23]_i_1_n_0 ),
        .Q(read_input[23]),
        .R(1'b0));
  FDRE \read_input_reg[24]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[24]_i_1_n_0 ),
        .Q(read_input[24]),
        .R(1'b0));
  FDRE \read_input_reg[25]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[25]_i_1_n_0 ),
        .Q(read_input[25]),
        .R(1'b0));
  FDRE \read_input_reg[26]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[26]_i_1_n_0 ),
        .Q(read_input[26]),
        .R(1'b0));
  FDRE \read_input_reg[27]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[27]_i_1_n_0 ),
        .Q(read_input[27]),
        .R(1'b0));
  FDRE \read_input_reg[28]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[28]_i_1_n_0 ),
        .Q(read_input[28]),
        .R(1'b0));
  FDRE \read_input_reg[29]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[29]_i_1_n_0 ),
        .Q(read_input[29]),
        .R(1'b0));
  FDRE \read_input_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[2]_i_1_n_0 ),
        .Q(read_input[2]),
        .R(1'b0));
  FDRE \read_input_reg[30]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[30]_i_1_n_0 ),
        .Q(read_input[30]),
        .R(1'b0));
  FDRE \read_input_reg[31]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[31]_i_2_n_0 ),
        .Q(read_input[31]),
        .R(1'b0));
  FDRE \read_input_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[3]_i_1_n_0 ),
        .Q(read_input[3]),
        .R(1'b0));
  FDRE \read_input_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[4]_i_1_n_0 ),
        .Q(read_input[4]),
        .R(1'b0));
  FDRE \read_input_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[5]_i_1_n_0 ),
        .Q(read_input[5]),
        .R(1'b0));
  FDRE \read_input_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[6]_i_1_n_0 ),
        .Q(read_input[6]),
        .R(1'b0));
  FDRE \read_input_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[7]_i_1_n_0 ),
        .Q(read_input[7]),
        .R(1'b0));
  FDRE \read_input_reg[8]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[8]_i_1_n_0 ),
        .Q(read_input[8]),
        .R(1'b0));
  FDRE \read_input_reg[9]
       (.C(ETH_CLK_OBUF),
        .CE(\read_input[31]_i_1_n_0 ),
        .D(\write_output[9]_i_1_n_0 ),
        .Q(read_input[9]),
        .R(1'b0));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_UNIQ_BASE_ registers_reg_r1_0_15_0_5
       (.ADDRA({1'b0,address_b_2}),
        .ADDRB({1'b0,address_b_2}),
        .ADDRC({1'b0,address_b_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[1:0]),
        .DIB(result[3:2]),
        .DIC(result[5:4]),
        .DID({1'b0,1'b0}),
        .DOA(register_b[1:0]),
        .DOB(register_b[3:2]),
        .DOC(register_b[5:4]),
        .DOD(NLW_registers_reg_r1_0_15_0_5_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD5 registers_reg_r1_0_15_12_17
       (.ADDRA({1'b0,address_b_2}),
        .ADDRB({1'b0,address_b_2}),
        .ADDRC({1'b0,address_b_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[13:12]),
        .DIB(result[15:14]),
        .DIC(result[17:16]),
        .DID({1'b0,1'b0}),
        .DOA(register_b[13:12]),
        .DOB(register_b[15:14]),
        .DOC(register_b[17:16]),
        .DOD(NLW_registers_reg_r1_0_15_12_17_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD6 registers_reg_r1_0_15_18_23
       (.ADDRA({1'b0,address_b_2}),
        .ADDRB({1'b0,address_b_2}),
        .ADDRC({1'b0,address_b_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[19:18]),
        .DIB(result[21:20]),
        .DIC(result[23:22]),
        .DID({1'b0,1'b0}),
        .DOA(register_b[19:18]),
        .DOB(register_b[21:20]),
        .DOC(register_b[23:22]),
        .DOD(NLW_registers_reg_r1_0_15_18_23_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD7 registers_reg_r1_0_15_24_29
       (.ADDRA({1'b0,address_b_2}),
        .ADDRB({1'b0,address_b_2}),
        .ADDRC({1'b0,address_b_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[25:24]),
        .DIB(result[27:26]),
        .DIC(result[29:28]),
        .DID({1'b0,1'b0}),
        .DOA(register_b[25:24]),
        .DOB(register_b[27:26]),
        .DOC(register_b[29:28]),
        .DOD(NLW_registers_reg_r1_0_15_24_29_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD8 registers_reg_r1_0_15_30_31
       (.ADDRA({1'b0,address_b_2}),
        .ADDRB({1'b0,address_b_2}),
        .ADDRC({1'b0,address_b_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[31:30]),
        .DIB({1'b0,1'b0}),
        .DIC({1'b0,1'b0}),
        .DID({1'b0,1'b0}),
        .DOA(register_b[31:30]),
        .DOB(NLW_registers_reg_r1_0_15_30_31_DOB_UNCONNECTED[1:0]),
        .DOC(NLW_registers_reg_r1_0_15_30_31_DOC_UNCONNECTED[1:0]),
        .DOD(NLW_registers_reg_r1_0_15_30_31_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD4 registers_reg_r1_0_15_6_11
       (.ADDRA({1'b0,address_b_2}),
        .ADDRB({1'b0,address_b_2}),
        .ADDRC({1'b0,address_b_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[7:6]),
        .DIB(result[9:8]),
        .DIC(result[11:10]),
        .DID({1'b0,1'b0}),
        .DOA(register_b[7:6]),
        .DOB(register_b[9:8]),
        .DOC(register_b[11:10]),
        .DOD(NLW_registers_reg_r1_0_15_6_11_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD9 registers_reg_r2_0_15_0_5
       (.ADDRA({1'b0,address_a_2}),
        .ADDRB({1'b0,address_a_2}),
        .ADDRC({1'b0,address_a_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[1:0]),
        .DIB(result[3:2]),
        .DIC(result[5:4]),
        .DID({1'b0,1'b0}),
        .DOA(register_a[1:0]),
        .DOB(register_a[3:2]),
        .DOC(register_a[5:4]),
        .DOD(NLW_registers_reg_r2_0_15_0_5_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD11 registers_reg_r2_0_15_12_17
       (.ADDRA({1'b0,address_a_2}),
        .ADDRB({1'b0,address_a_2}),
        .ADDRC({1'b0,address_a_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[13:12]),
        .DIB(result[15:14]),
        .DIC(result[17:16]),
        .DID({1'b0,1'b0}),
        .DOA(register_a[13:12]),
        .DOB(register_a[15:14]),
        .DOC(register_a[17:16]),
        .DOD(NLW_registers_reg_r2_0_15_12_17_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD12 registers_reg_r2_0_15_18_23
       (.ADDRA({1'b0,address_a_2}),
        .ADDRB({1'b0,address_a_2}),
        .ADDRC({1'b0,address_a_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[19:18]),
        .DIB(result[21:20]),
        .DIC(result[23:22]),
        .DID({1'b0,1'b0}),
        .DOA(register_a[19:18]),
        .DOB(register_a[21:20]),
        .DOC(register_a[23:22]),
        .DOD(NLW_registers_reg_r2_0_15_18_23_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD13 registers_reg_r2_0_15_24_29
       (.ADDRA({1'b0,address_a_2}),
        .ADDRB({1'b0,address_a_2}),
        .ADDRC({1'b0,address_a_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[25:24]),
        .DIB(result[27:26]),
        .DIC(result[29:28]),
        .DID({1'b0,1'b0}),
        .DOA(register_a[25:24]),
        .DOB(register_a[27:26]),
        .DOC(register_a[29:28]),
        .DOD(NLW_registers_reg_r2_0_15_24_29_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD14 registers_reg_r2_0_15_30_31
       (.ADDRA({1'b0,address_a_2}),
        .ADDRB({1'b0,address_a_2}),
        .ADDRC({1'b0,address_a_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[31:30]),
        .DIB({1'b0,1'b0}),
        .DIC({1'b0,1'b0}),
        .DID({1'b0,1'b0}),
        .DOA(register_a[31:30]),
        .DOB(NLW_registers_reg_r2_0_15_30_31_DOB_UNCONNECTED[1:0]),
        .DOC(NLW_registers_reg_r2_0_15_30_31_DOC_UNCONNECTED[1:0]),
        .DOD(NLW_registers_reg_r2_0_15_30_31_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  (* INIT_A = "64'h0000000000000000" *)
  (* INIT_B = "64'h0000000000000000" *)
  (* INIT_C = "64'h0000000000000000" *)
  (* INIT_D = "64'h0000000000000000" *)
  RAM32M_HD10 registers_reg_r2_0_15_6_11
       (.ADDRA({1'b0,address_a_2}),
        .ADDRB({1'b0,address_a_2}),
        .ADDRC({1'b0,address_a_2}),
        .ADDRD({1'b0,address_z_3}),
        .DIA(result[7:6]),
        .DIB(result[9:8]),
        .DIC(result[11:10]),
        .DID({1'b0,1'b0}),
        .DOA(register_a[7:6]),
        .DOB(register_a[9:8]),
        .DOC(register_a[11:10]),
        .DOD(NLW_registers_reg_r2_0_15_6_11_DOD_UNCONNECTED[1:0]),
        .WCLK(ETH_CLK_OBUF),
        .WE(write_enable));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[0]_i_1
       (.I0(\result[0]_i_2_n_0 ),
        .I1(\result_reg[3]_i_3_n_7 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result[0]_i_3_n_0 ),
        .I4(\result[7]_i_5_n_0 ),
        .I5(data5[0]),
        .O(\result[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_10
       (.I0(\write_output[24]_i_1_n_0 ),
        .I1(store_data[26]),
        .I2(store_data[24]),
        .I3(store_data[25]),
        .I4(\write_output[26]_i_1_n_0 ),
        .I5(\write_output[25]_i_1_n_0 ),
        .O(\result[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_12
       (.I0(\write_output[21]_i_1_n_0 ),
        .I1(store_data[23]),
        .I2(store_data[21]),
        .I3(store_data[22]),
        .I4(\write_output[23]_i_1_n_0 ),
        .I5(\write_output[22]_i_1_n_0 ),
        .O(\result[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_13
       (.I0(\write_output[18]_i_1_n_0 ),
        .I1(store_data[20]),
        .I2(store_data[18]),
        .I3(store_data[19]),
        .I4(\write_output[20]_i_1_n_0 ),
        .I5(\write_output[19]_i_1_n_0 ),
        .O(\result[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_14
       (.I0(\write_output[15]_i_1_n_0 ),
        .I1(store_data[17]),
        .I2(store_data[15]),
        .I3(store_data[16]),
        .I4(\write_output[17]_i_1_n_0 ),
        .I5(\write_output[16]_i_1_n_0 ),
        .O(\result[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_15
       (.I0(\write_output[12]_i_1_n_0 ),
        .I1(store_data[14]),
        .I2(store_data[12]),
        .I3(store_data[13]),
        .I4(\write_output[14]_i_1_n_0 ),
        .I5(\write_output[13]_i_1_n_0 ),
        .O(\result[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_16
       (.I0(\write_output[9]_i_1_n_0 ),
        .I1(store_data[11]),
        .I2(store_data[9]),
        .I3(store_data[10]),
        .I4(\write_output[11]_i_1_n_0 ),
        .I5(\write_output[10]_i_1_n_0 ),
        .O(\result[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_17
       (.I0(\write_output[6]_i_1_n_0 ),
        .I1(store_data[8]),
        .I2(store_data[6]),
        .I3(store_data[7]),
        .I4(\write_output[8]_i_1_n_0 ),
        .I5(\write_output[7]_i_1_n_0 ),
        .O(\result[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_18
       (.I0(\write_output[3]_i_1_n_0 ),
        .I1(store_data[5]),
        .I2(store_data[3]),
        .I3(store_data[4]),
        .I4(\write_output[5]_i_1_n_0 ),
        .I5(\write_output[4]_i_1_n_0 ),
        .O(\result[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_19
       (.I0(\write_output[0]_i_1_n_0 ),
        .I1(store_data[2]),
        .I2(store_data[0]),
        .I3(store_data[1]),
        .I4(\write_output[2]_i_1_n_0 ),
        .I5(\write_output[1]_i_1_n_0 ),
        .O(\result[0]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4000))
    \result[0]_i_2
       (.I0(opcode_2[3]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[2]),
        .I3(\result_reg[0]_i_4_n_1 ),
        .I4(\result[0]_i_5_n_0 ),
        .O(\result[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAEABAFAAAEAAAEA))
    \result[0]_i_3
       (.I0(\result[0]_i_6_n_0 ),
        .I1(opcode_2[1]),
        .I2(memory_reg_0_i_2_n_0),
        .I3(program_counter_2[0]),
        .I4(opcode_2[0]),
        .I5(address_b_2[0]),
        .O(\result[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00F0444400004444))
    \result[0]_i_5
       (.I0(\state_reg_n_0_[1] ),
        .I1(load_data[0]),
        .I2(data4[0]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[3]),
        .O(\result[0]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h0C000A00))
    \result[0]_i_6
       (.I0(DATA[0]),
        .I1(OUT1[0]),
        .I2(\state_reg_n_0_[0] ),
        .I3(\state_reg_n_0_[1] ),
        .I4(read_input[1]),
        .O(\result[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hE2001D0000E2001D))
    \result[0]_i_8
       (.I0(register_a[31]),
        .I1(operand_a1),
        .I2(result[31]),
        .I3(\write_output[30]_i_1_n_0 ),
        .I4(store_data[31]),
        .I5(store_data[30]),
        .O(\result[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h8400210000840021))
    \result[0]_i_9
       (.I0(\write_output[27]_i_1_n_0 ),
        .I1(store_data[29]),
        .I2(store_data[27]),
        .I3(store_data[28]),
        .I4(\write_output[29]_i_1_n_0 ),
        .I5(\write_output[28]_i_1_n_0 ),
        .O(\result[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFAEFFAEFFAE))
    \result[10]_i_1
       (.I0(\result[10]_i_2_n_0 ),
        .I1(load_data[10]),
        .I2(\result[11]_i_3_n_0 ),
        .I3(\result[31]_i_7_n_0 ),
        .I4(\result[16]_i_5_n_0 ),
        .I5(data4[10]),
        .O(\result[10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \result[10]_i_2
       (.I0(\result_reg[11]_i_5_n_5 ),
        .I1(\result[16]_i_3_n_0 ),
        .I2(\result[7]_i_5_n_0 ),
        .I3(data5[10]),
        .I4(\result[16]_i_7_n_0 ),
        .I5(data2[10]),
        .O(\result[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFAEFFAEFFAE))
    \result[11]_i_1
       (.I0(\result[11]_i_2_n_0 ),
        .I1(load_data[11]),
        .I2(\result[11]_i_3_n_0 ),
        .I3(\result[31]_i_7_n_0 ),
        .I4(\result[16]_i_5_n_0 ),
        .I5(data4[11]),
        .O(\result[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[11]_i_10
       (.I0(register_a[8]),
        .I1(operand_a1),
        .I2(register_b[8]),
        .I3(operand_b1),
        .I4(result[8]),
        .O(\result[11]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[11]_i_11
       (.I0(register_a[11]),
        .I1(operand_a1),
        .I2(result[11]),
        .I3(literal_2[15]),
        .O(\result[11]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[11]_i_12
       (.I0(register_a[10]),
        .I1(operand_a1),
        .I2(result[10]),
        .I3(literal_2[15]),
        .O(\result[11]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[11]_i_13
       (.I0(register_a[9]),
        .I1(operand_a1),
        .I2(result[9]),
        .I3(literal_2[9]),
        .O(\result[11]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[11]_i_14
       (.I0(register_a[8]),
        .I1(operand_a1),
        .I2(result[8]),
        .I3(literal_2[8]),
        .O(\result[11]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[11]_i_15
       (.I0(result[7]),
        .I1(operand_b1),
        .I2(register_b[7]),
        .I3(operand_a1),
        .I4(register_a[7]),
        .O(\result[11]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[11]_i_16
       (.I0(result[6]),
        .I1(operand_b1),
        .I2(register_b[6]),
        .I3(operand_a1),
        .I4(register_a[6]),
        .O(\result[11]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[11]_i_17
       (.I0(result[5]),
        .I1(operand_b1),
        .I2(register_b[5]),
        .I3(operand_a1),
        .I4(register_a[5]),
        .O(\result[11]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[11]_i_18
       (.I0(result[4]),
        .I1(operand_b1),
        .I2(register_b[4]),
        .I3(operand_a1),
        .I4(register_a[4]),
        .O(\result[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888))
    \result[11]_i_2
       (.I0(\result_reg[11]_i_5_n_4 ),
        .I1(\result[16]_i_3_n_0 ),
        .I2(\result[7]_i_5_n_0 ),
        .I3(data5[11]),
        .I4(\result[16]_i_7_n_0 ),
        .I5(data2[11]),
        .O(\result[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE))
    \result[11]_i_3
       (.I0(\state_reg_n_0_[0] ),
        .I1(\state_reg_n_0_[1] ),
        .O(\result[11]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[11]_i_7
       (.I0(register_a[11]),
        .I1(operand_a1),
        .I2(register_b[11]),
        .I3(operand_b1),
        .I4(result[11]),
        .O(\result[11]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[11]_i_8
       (.I0(register_a[10]),
        .I1(operand_a1),
        .I2(register_b[10]),
        .I3(operand_b1),
        .I4(result[10]),
        .O(\result[11]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[11]_i_9
       (.I0(register_a[9]),
        .I1(operand_a1),
        .I2(register_b[9]),
        .I3(operand_b1),
        .I4(result[9]),
        .O(\result[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAAAAA))
    \result[12]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[2]),
        .I4(data4[12]),
        .I5(\result[12]_i_2_n_0 ),
        .O(\result[12]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF020202))
    \result[12]_i_2
       (.I0(load_data[12]),
        .I1(\state_reg_n_0_[1] ),
        .I2(\state_reg_n_0_[0] ),
        .I3(\result[16]_i_7_n_0 ),
        .I4(data2[12]),
        .I5(\result[12]_i_4_n_0 ),
        .O(\result[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF888888888888888))
    \result[12]_i_4
       (.I0(\result[16]_i_3_n_0 ),
        .I1(\result_reg[16]_i_9_n_7 ),
        .I2(data5[12]),
        .I3(opcode_2[3]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[2]),
        .O(\result[12]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAAAAA))
    \result[13]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[2]),
        .I4(data4[13]),
        .I5(\result[13]_i_2_n_0 ),
        .O(\result[13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8))
    \result[13]_i_2
       (.I0(\result[16]_i_7_n_0 ),
        .I1(data2[13]),
        .I2(load_data[13]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\state_reg_n_0_[0] ),
        .I5(\result[13]_i_3_n_0 ),
        .O(\result[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF800080008000))
    \result[13]_i_3
       (.I0(data5[13]),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[2]),
        .I4(\result_reg[16]_i_9_n_6 ),
        .I5(\result[16]_i_3_n_0 ),
        .O(\result[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAAAAA))
    \result[14]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[2]),
        .I4(data4[14]),
        .I5(\result[14]_i_2_n_0 ),
        .O(\result[14]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8))
    \result[14]_i_2
       (.I0(\result[16]_i_7_n_0 ),
        .I1(data2[14]),
        .I2(load_data[14]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\state_reg_n_0_[0] ),
        .I5(\result[14]_i_3_n_0 ),
        .O(\result[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF800080008000))
    \result[14]_i_3
       (.I0(data5[14]),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[2]),
        .I4(\result_reg[16]_i_9_n_5 ),
        .I5(\result[16]_i_3_n_0 ),
        .O(\result[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAAAAA))
    \result[15]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[2]),
        .I4(data4[15]),
        .I5(\result[15]_i_3_n_0 ),
        .O(\result[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888F8))
    \result[15]_i_3
       (.I0(\result[16]_i_7_n_0 ),
        .I1(data2[15]),
        .I2(load_data[15]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\state_reg_n_0_[0] ),
        .I5(\result[15]_i_8_n_0 ),
        .O(\result[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[15]_i_4
       (.I0(result[15]),
        .I1(operand_b1),
        .I2(register_b[15]),
        .I3(operand_a1),
        .I4(register_a[15]),
        .O(\result[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[15]_i_5
       (.I0(result[14]),
        .I1(operand_b1),
        .I2(register_b[14]),
        .I3(operand_a1),
        .I4(register_a[14]),
        .O(\result[15]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[15]_i_6
       (.I0(result[13]),
        .I1(operand_b1),
        .I2(register_b[13]),
        .I3(operand_a1),
        .I4(register_a[13]),
        .O(\result[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[15]_i_7
       (.I0(result[12]),
        .I1(operand_b1),
        .I2(register_b[12]),
        .I3(operand_a1),
        .I4(register_a[12]),
        .O(\result[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF800080008000))
    \result[15]_i_8
       (.I0(data5[15]),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[2]),
        .I4(\result_reg[16]_i_9_n_4 ),
        .I5(\result[16]_i_3_n_0 ),
        .O(\result[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[16]_i_1
       (.I0(\result[16]_i_2_n_0 ),
        .I1(\result[16]_i_3_n_0 ),
        .I2(\result_reg[16]_i_4_n_7 ),
        .I3(\result[31]_i_7_n_0 ),
        .I4(\result[16]_i_5_n_0 ),
        .I5(data4[16]),
        .O(\result[16]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[16]_i_10
       (.I0(result[19]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[19]),
        .O(\result[16]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[16]_i_11
       (.I0(result[18]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[18]),
        .O(\result[16]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[16]_i_12
       (.I0(result[17]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[17]),
        .O(\result[16]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[16]_i_13
       (.I0(result[16]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[16]),
        .O(\result[16]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[16]_i_14
       (.I0(register_a[19]),
        .I1(operand_a1),
        .I2(register_b[19]),
        .I3(operand_b1),
        .I4(result[19]),
        .O(\result[16]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[16]_i_15
       (.I0(register_a[18]),
        .I1(operand_a1),
        .I2(register_b[18]),
        .I3(operand_b1),
        .I4(result[18]),
        .O(\result[16]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[16]_i_16
       (.I0(register_a[17]),
        .I1(operand_a1),
        .I2(register_b[17]),
        .I3(operand_b1),
        .I4(result[17]),
        .O(\result[16]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[16]_i_17
       (.I0(register_a[16]),
        .I1(operand_a1),
        .I2(register_b[16]),
        .I3(operand_b1),
        .I4(result[16]),
        .O(\result[16]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[16]_i_2
       (.I0(data5[16]),
        .I1(\result[7]_i_5_n_0 ),
        .I2(\result[16]_i_7_n_0 ),
        .I3(data2[16]),
        .I4(load_data[16]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[16]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[16]_i_21
       (.I0(register_a[15]),
        .I1(operand_a1),
        .I2(result[15]),
        .I3(literal_2[15]),
        .O(\result[16]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[16]_i_22
       (.I0(register_a[14]),
        .I1(operand_a1),
        .I2(result[14]),
        .I3(literal_2[15]),
        .O(\result[16]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[16]_i_23
       (.I0(register_a[13]),
        .I1(operand_a1),
        .I2(result[13]),
        .I3(literal_2[15]),
        .O(\result[16]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[16]_i_24
       (.I0(register_a[12]),
        .I1(operand_a1),
        .I2(result[12]),
        .I3(literal_2[15]),
        .O(\result[16]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h00000400))
    \result[16]_i_3
       (.I0(opcode_2[3]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[2]),
        .I3(opcode_2[0]),
        .I4(opcode_2[1]),
        .O(\result[16]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h40))
    \result[16]_i_5
       (.I0(opcode_2[2]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[3]),
        .O(\result[16]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0400))
    \result[16]_i_7
       (.I0(opcode_2[3]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[2]),
        .I3(opcode_2[1]),
        .O(\result[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[17]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[17]),
        .I5(\result[17]_i_2_n_0 ),
        .O(\result[17]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[17]_i_2
       (.I0(data4[17]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[16]_i_4_n_6 ),
        .I4(load_data[17]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[18]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[18]),
        .I5(\result[18]_i_2_n_0 ),
        .O(\result[18]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[18]_i_2
       (.I0(data4[18]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[16]_i_4_n_5 ),
        .I4(load_data[18]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[19]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[19]),
        .I5(\result[19]_i_3_n_0 ),
        .O(\result[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[19]_i_10
       (.I0(register_a[14]),
        .I1(operand_a1),
        .I2(register_b[14]),
        .I3(operand_b1),
        .I4(result[14]),
        .O(\result[19]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[19]_i_11
       (.I0(register_a[13]),
        .I1(operand_a1),
        .I2(register_b[13]),
        .I3(operand_b1),
        .I4(result[13]),
        .O(\result[19]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[19]_i_12
       (.I0(register_a[12]),
        .I1(operand_a1),
        .I2(register_b[12]),
        .I3(operand_b1),
        .I4(result[12]),
        .O(\result[19]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[19]_i_3
       (.I0(data4[19]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[16]_i_4_n_4 ),
        .I4(load_data[19]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[19]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[19]_i_5
       (.I0(result[19]),
        .I1(operand_b1),
        .I2(register_b[19]),
        .I3(operand_a1),
        .I4(register_a[19]),
        .O(\result[19]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[19]_i_6
       (.I0(result[18]),
        .I1(operand_b1),
        .I2(register_b[18]),
        .I3(operand_a1),
        .I4(register_a[18]),
        .O(\result[19]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[19]_i_7
       (.I0(result[17]),
        .I1(operand_b1),
        .I2(register_b[17]),
        .I3(operand_a1),
        .I4(register_a[17]),
        .O(\result[19]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[19]_i_8
       (.I0(result[16]),
        .I1(operand_b1),
        .I2(register_b[16]),
        .I3(operand_a1),
        .I4(register_a[16]),
        .O(\result[19]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[19]_i_9
       (.I0(register_a[15]),
        .I1(operand_a1),
        .I2(register_b[15]),
        .I3(operand_b1),
        .I4(result[15]),
        .O(\result[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[1]_i_1
       (.I0(\result[1]_i_2_n_0 ),
        .I1(\result_reg[3]_i_3_n_6 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result[1]_i_3_n_0 ),
        .I4(\result[7]_i_5_n_0 ),
        .I5(data5[1]),
        .O(\result[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00F0444400004444))
    \result[1]_i_2
       (.I0(\state_reg_n_0_[1] ),
        .I1(load_data[1]),
        .I2(data4[1]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[3]),
        .O(\result[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEECFCCCCEECCCCCC))
    \result[1]_i_3
       (.I0(data2[1]),
        .I1(\result[1]_i_4_n_0 ),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(memory_reg_0_i_2_n_0),
        .I5(address_b_2[1]),
        .O(\result[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0C000A00))
    \result[1]_i_4
       (.I0(DATA[1]),
        .I1(OUT1[1]),
        .I2(\state_reg_n_0_[0] ),
        .I3(\state_reg_n_0_[1] ),
        .I4(read_input[1]),
        .O(\result[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[20]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[20]),
        .I5(\result[20]_i_2_n_0 ),
        .O(\result[20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[20]_i_2
       (.I0(data4[20]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[23]_i_9_n_7 ),
        .I4(load_data[20]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[21]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[21]),
        .I5(\result[21]_i_2_n_0 ),
        .O(\result[21]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[21]_i_2
       (.I0(data4[21]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[23]_i_9_n_6 ),
        .I4(load_data[21]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[22]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[22]),
        .I5(\result[22]_i_2_n_0 ),
        .O(\result[22]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[22]_i_2
       (.I0(data4[22]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[23]_i_9_n_5 ),
        .I4(load_data[22]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[22]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[23]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[23]),
        .I5(\result[23]_i_3_n_0 ),
        .O(\result[23]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[23]_i_10
       (.I0(register_a[23]),
        .I1(operand_a1),
        .I2(register_b[23]),
        .I3(operand_b1),
        .I4(result[23]),
        .O(\result[23]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[23]_i_11
       (.I0(register_a[22]),
        .I1(operand_a1),
        .I2(register_b[22]),
        .I3(operand_b1),
        .I4(result[22]),
        .O(\result[23]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[23]_i_12
       (.I0(register_a[21]),
        .I1(operand_a1),
        .I2(register_b[21]),
        .I3(operand_b1),
        .I4(result[21]),
        .O(\result[23]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[23]_i_13
       (.I0(register_a[20]),
        .I1(operand_a1),
        .I2(register_b[20]),
        .I3(operand_b1),
        .I4(result[20]),
        .O(\result[23]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[23]_i_14
       (.I0(result[23]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[23]),
        .O(\result[23]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[23]_i_15
       (.I0(result[22]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[22]),
        .O(\result[23]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[23]_i_16
       (.I0(result[21]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[21]),
        .O(\result[23]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[23]_i_17
       (.I0(result[20]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[20]),
        .O(\result[23]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[23]_i_3
       (.I0(data4[23]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[23]_i_9_n_4 ),
        .I4(load_data[23]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[23]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[23]_i_4
       (.I0(result[23]),
        .I1(operand_b1),
        .I2(register_b[23]),
        .I3(operand_a1),
        .I4(register_a[23]),
        .O(\result[23]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[23]_i_5
       (.I0(result[22]),
        .I1(operand_b1),
        .I2(register_b[22]),
        .I3(operand_a1),
        .I4(register_a[22]),
        .O(\result[23]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[23]_i_6
       (.I0(result[21]),
        .I1(operand_b1),
        .I2(register_b[21]),
        .I3(operand_a1),
        .I4(register_a[21]),
        .O(\result[23]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[23]_i_7
       (.I0(result[20]),
        .I1(operand_b1),
        .I2(register_b[20]),
        .I3(operand_a1),
        .I4(register_a[20]),
        .O(\result[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[24]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[24]),
        .I5(\result[24]_i_2_n_0 ),
        .O(\result[24]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[24]_i_2
       (.I0(data4[24]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[27]_i_9_n_7 ),
        .I4(load_data[24]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[24]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[25]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[25]),
        .I5(\result[25]_i_2_n_0 ),
        .O(\result[25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[25]_i_2
       (.I0(data4[25]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[27]_i_9_n_6 ),
        .I4(load_data[25]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[25]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[26]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[26]),
        .I5(\result[26]_i_2_n_0 ),
        .O(\result[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[26]_i_2
       (.I0(data4[26]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[27]_i_9_n_5 ),
        .I4(load_data[26]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[26]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[27]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[27]),
        .I5(\result[27]_i_3_n_0 ),
        .O(\result[27]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[27]_i_10
       (.I0(register_a[27]),
        .I1(operand_a1),
        .I2(register_b[27]),
        .I3(operand_b1),
        .I4(result[27]),
        .O(\result[27]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[27]_i_11
       (.I0(register_a[26]),
        .I1(operand_a1),
        .I2(register_b[26]),
        .I3(operand_b1),
        .I4(result[26]),
        .O(\result[27]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[27]_i_12
       (.I0(register_a[25]),
        .I1(operand_a1),
        .I2(register_b[25]),
        .I3(operand_b1),
        .I4(result[25]),
        .O(\result[27]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[27]_i_13
       (.I0(register_a[24]),
        .I1(operand_a1),
        .I2(register_b[24]),
        .I3(operand_b1),
        .I4(result[24]),
        .O(\result[27]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[27]_i_14
       (.I0(result[27]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[27]),
        .O(\result[27]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[27]_i_15
       (.I0(result[26]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[26]),
        .O(\result[27]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[27]_i_16
       (.I0(result[25]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[25]),
        .O(\result[27]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[27]_i_17
       (.I0(result[24]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[24]),
        .O(\result[27]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[27]_i_3
       (.I0(data4[27]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[27]_i_9_n_4 ),
        .I4(load_data[27]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[27]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[27]_i_4
       (.I0(result[27]),
        .I1(operand_a1),
        .I2(register_a[27]),
        .I3(operand_b1),
        .I4(register_b[27]),
        .O(\result[27]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[27]_i_5
       (.I0(result[26]),
        .I1(operand_a1),
        .I2(register_a[26]),
        .I3(operand_b1),
        .I4(register_b[26]),
        .O(\result[27]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[27]_i_6
       (.I0(result[25]),
        .I1(operand_b1),
        .I2(register_b[25]),
        .I3(operand_a1),
        .I4(register_a[25]),
        .O(\result[27]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[27]_i_7
       (.I0(result[24]),
        .I1(operand_a1),
        .I2(register_a[24]),
        .I3(operand_b1),
        .I4(register_b[24]),
        .O(\result[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[28]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[28]),
        .I5(\result[28]_i_2_n_0 ),
        .O(\result[28]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[28]_i_2
       (.I0(data4[28]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[31]_i_17_n_7 ),
        .I4(load_data[28]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[28]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[29]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[29]),
        .I5(\result[29]_i_2_n_0 ),
        .O(\result[29]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[29]_i_2
       (.I0(data4[29]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[31]_i_17_n_6 ),
        .I4(load_data[29]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[29]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[2]_i_1
       (.I0(\result[2]_i_2_n_0 ),
        .I1(\result_reg[3]_i_3_n_5 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result[2]_i_3_n_0 ),
        .I4(\result[7]_i_5_n_0 ),
        .I5(data5[2]),
        .O(\result[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00F0444400004444))
    \result[2]_i_2
       (.I0(\state_reg_n_0_[1] ),
        .I1(load_data[2]),
        .I2(data4[2]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[3]),
        .O(\result[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEECFCCCCEECCCCCC))
    \result[2]_i_3
       (.I0(data2[2]),
        .I1(\result[2]_i_4_n_0 ),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(memory_reg_0_i_2_n_0),
        .I5(address_b_2[2]),
        .O(\result[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0C000A00))
    \result[2]_i_4
       (.I0(DATA[2]),
        .I1(OUT1[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(\state_reg_n_0_[1] ),
        .I4(read_input[1]),
        .O(\result[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[30]_i_1
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[30]),
        .I5(\result[30]_i_2_n_0 ),
        .O(\result[30]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[30]_i_2
       (.I0(data4[30]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[31]_i_17_n_5 ),
        .I4(load_data[30]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF02000222))
    \result[31]_i_1
       (.I0(\result[31]_i_3_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(OUT1_STB_reg),
        .I3(read_input[1]),
        .I4(S_DATA_STB_reg),
        .I5(\result[31]_i_6_n_0 ),
        .O(\result[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000))
    \result[31]_i_10
       (.I0(\result[31]_i_18_n_0 ),
        .I1(\result[31]_i_19_n_0 ),
        .I2(\result[31]_i_20_n_0 ),
        .I3(read_input[9]),
        .I4(\result[31]_i_21_n_0 ),
        .I5(\result[31]_i_22_n_0 ),
        .O(\result[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h1080000080800000))
    \result[31]_i_11
       (.I0(opcode_2[0]),
        .I1(opcode_2[1]),
        .I2(\state_reg_n_0_[1] ),
        .I3(opcode_2[3]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[2]),
        .O(\result[31]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[31]_i_12
       (.I0(result[31]),
        .I1(operand_a1),
        .I2(register_a[31]),
        .I3(operand_b1),
        .I4(register_b[31]),
        .O(\result[31]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[31]_i_13
       (.I0(result[30]),
        .I1(operand_b1),
        .I2(register_b[30]),
        .I3(operand_a1),
        .I4(register_a[30]),
        .O(\result[31]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[31]_i_14
       (.I0(result[29]),
        .I1(operand_a1),
        .I2(register_a[29]),
        .I3(operand_b1),
        .I4(register_b[29]),
        .O(\result[31]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[31]_i_15
       (.I0(result[28]),
        .I1(operand_b1),
        .I2(register_b[28]),
        .I3(operand_a1),
        .I4(register_a[28]),
        .O(\result[31]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001))
    \result[31]_i_18
       (.I0(read_input[7]),
        .I1(read_input[10]),
        .I2(read_input[14]),
        .I3(read_input[11]),
        .I4(read_input[8]),
        .I5(read_input[13]),
        .O(\result[31]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001))
    \result[31]_i_19
       (.I0(read_input[16]),
        .I1(read_input[15]),
        .I2(read_input[19]),
        .I3(read_input[20]),
        .I4(read_input[21]),
        .I5(read_input[22]),
        .O(\result[31]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA))
    \result[31]_i_2
       (.I0(\result[31]_i_7_n_0 ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[0] ),
        .I3(opcode_2[3]),
        .I4(data5[31]),
        .I5(\result[31]_i_9_n_0 ),
        .O(\result[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001))
    \result[31]_i_20
       (.I0(read_input[30]),
        .I1(read_input[29]),
        .I2(read_input[17]),
        .I3(read_input[18]),
        .I4(read_input[27]),
        .I5(read_input[28]),
        .O(\result[31]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001))
    \result[31]_i_21
       (.I0(read_input[4]),
        .I1(read_input[3]),
        .I2(read_input[23]),
        .I3(read_input[24]),
        .I4(read_input[25]),
        .I5(read_input[26]),
        .O(\result[31]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001))
    \result[31]_i_22
       (.I0(read_input[0]),
        .I1(read_input[12]),
        .I2(read_input[5]),
        .I3(read_input[6]),
        .I4(read_input[2]),
        .I5(read_input[31]),
        .O(\result[31]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h8008))
    \result[31]_i_23
       (.I0(\write_output[31]_i_4_n_0 ),
        .I1(write_enable),
        .I2(address_a_2[3]),
        .I3(address_z_3[3]),
        .O(operand_a1));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[31]_i_24
       (.I0(register_a[31]),
        .I1(operand_a1),
        .I2(register_b[31]),
        .I3(operand_b1),
        .I4(result[31]),
        .O(\result[31]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[31]_i_25
       (.I0(register_a[30]),
        .I1(operand_a1),
        .I2(register_b[30]),
        .I3(operand_b1),
        .I4(result[30]),
        .O(\result[31]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[31]_i_26
       (.I0(register_a[29]),
        .I1(operand_a1),
        .I2(register_b[29]),
        .I3(operand_b1),
        .I4(result[29]),
        .O(\result[31]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hEEE1DD2D))
    \result[31]_i_27
       (.I0(register_a[28]),
        .I1(operand_a1),
        .I2(register_b[28]),
        .I3(operand_b1),
        .I4(result[28]),
        .O(\result[31]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[31]_i_28
       (.I0(result[31]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[31]),
        .O(\result[31]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[31]_i_29
       (.I0(result[30]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[30]),
        .O(\result[31]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h8))
    \result[31]_i_3
       (.I0(\result[31]_i_10_n_0 ),
        .I1(\state_reg_n_0_[2] ),
        .O(\result[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[31]_i_30
       (.I0(result[29]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[29]),
        .O(\result[31]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \result[31]_i_31
       (.I0(result[28]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[28]),
        .O(\result[31]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h00F200F200F0FFF0))
    \result[31]_i_6
       (.I0(memory_reg_0_i_2_n_0),
        .I1(opcode_2[1]),
        .I2(\result[31]_i_11_n_0 ),
        .I3(\state_reg_n_0_[2] ),
        .I4(\state_reg_n_0_[0] ),
        .I5(\state_reg_n_0_[1] ),
        .O(\result[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000))
    \result[31]_i_7
       (.I0(opcode_2[0]),
        .I1(opcode_2[1]),
        .I2(opcode_2[2]),
        .I3(\state_reg_n_0_[0] ),
        .I4(opcode_2[3]),
        .I5(literal_2[15]),
        .O(\result[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF888F888FFFFF888))
    \result[31]_i_9
       (.I0(data4[31]),
        .I1(\result[16]_i_5_n_0 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result_reg[31]_i_17_n_4 ),
        .I4(load_data[31]),
        .I5(\result[11]_i_3_n_0 ),
        .O(\result[31]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[3]_i_1
       (.I0(\result[3]_i_2_n_0 ),
        .I1(\result_reg[3]_i_3_n_4 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result[3]_i_4_n_0 ),
        .I4(\result[7]_i_5_n_0 ),
        .I5(data5[3]),
        .O(\result[3]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[3]_i_10
       (.I0(register_a[0]),
        .I1(operand_a1),
        .I2(result[0]),
        .I3(address_b_2[0]),
        .O(\result[3]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h0C000A00))
    \result[3]_i_11
       (.I0(DATA[3]),
        .I1(OUT1[3]),
        .I2(\state_reg_n_0_[0] ),
        .I3(\state_reg_n_0_[1] ),
        .I4(read_input[1]),
        .O(\result[3]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[3]_i_12
       (.I0(register_a[3]),
        .I1(operand_a1),
        .I2(register_b[3]),
        .I3(operand_b1),
        .I4(result[3]),
        .O(\result[3]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[3]_i_13
       (.I0(register_a[2]),
        .I1(operand_a1),
        .I2(register_b[2]),
        .I3(operand_b1),
        .I4(result[2]),
        .O(\result[3]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[3]_i_14
       (.I0(register_a[1]),
        .I1(operand_a1),
        .I2(register_b[1]),
        .I3(operand_b1),
        .I4(result[1]),
        .O(\result[3]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[3]_i_15
       (.I0(register_a[0]),
        .I1(operand_a1),
        .I2(register_b[0]),
        .I3(operand_b1),
        .I4(result[0]),
        .O(\result[3]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[3]_i_16
       (.I0(result[3]),
        .I1(operand_b1),
        .I2(register_b[3]),
        .I3(operand_a1),
        .I4(register_a[3]),
        .O(\result[3]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[3]_i_17
       (.I0(result[2]),
        .I1(operand_b1),
        .I2(register_b[2]),
        .I3(operand_a1),
        .I4(register_a[2]),
        .O(\result[3]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[3]_i_18
       (.I0(result[1]),
        .I1(operand_b1),
        .I2(register_b[1]),
        .I3(operand_a1),
        .I4(register_a[1]),
        .O(\result[3]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hEDB8ED47))
    \result[3]_i_19
       (.I0(result[0]),
        .I1(operand_b1),
        .I2(register_b[0]),
        .I3(operand_a1),
        .I4(register_a[0]),
        .O(\result[3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00F0444400004444))
    \result[3]_i_2
       (.I0(\state_reg_n_0_[1] ),
        .I1(load_data[3]),
        .I2(data4[3]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[3]),
        .O(\result[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEECFCCCCEECCCCCC))
    \result[3]_i_4
       (.I0(data2[3]),
        .I1(\result[3]_i_11_n_0 ),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(memory_reg_0_i_2_n_0),
        .I5(address_b_2[3]),
        .O(\result[3]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[3]_i_7
       (.I0(register_a[3]),
        .I1(operand_a1),
        .I2(result[3]),
        .I3(address_b_2[3]),
        .O(\result[3]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[3]_i_8
       (.I0(register_a[2]),
        .I1(operand_a1),
        .I2(result[2]),
        .I3(address_b_2[2]),
        .O(\result[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[3]_i_9
       (.I0(register_a[1]),
        .I1(operand_a1),
        .I2(result[1]),
        .I3(address_b_2[1]),
        .O(\result[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[4]_i_1
       (.I0(\result[4]_i_2_n_0 ),
        .I1(\result_reg[7]_i_3_n_7 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result[4]_i_3_n_0 ),
        .I4(\result[7]_i_5_n_0 ),
        .I5(data5[4]),
        .O(\result[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00F0444400004444))
    \result[4]_i_2
       (.I0(\state_reg_n_0_[1] ),
        .I1(load_data[4]),
        .I2(data4[4]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[3]),
        .O(\result[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEECFCCCCEECCCCCC))
    \result[4]_i_3
       (.I0(data2[4]),
        .I1(\result[4]_i_5_n_0 ),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(memory_reg_0_i_2_n_0),
        .I5(literal_2[4]),
        .O(\result[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0C000A00))
    \result[4]_i_5
       (.I0(DATA[4]),
        .I1(OUT1[4]),
        .I2(\state_reg_n_0_[0] ),
        .I3(\state_reg_n_0_[1] ),
        .I4(read_input[1]),
        .O(\result[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[5]_i_1
       (.I0(\result[5]_i_2_n_0 ),
        .I1(\result_reg[7]_i_3_n_6 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result[5]_i_3_n_0 ),
        .I4(\result[7]_i_5_n_0 ),
        .I5(data5[5]),
        .O(\result[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00F0444400004444))
    \result[5]_i_2
       (.I0(\state_reg_n_0_[1] ),
        .I1(load_data[5]),
        .I2(data4[5]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[3]),
        .O(\result[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEECFCCCCEECCCCCC))
    \result[5]_i_3
       (.I0(data2[5]),
        .I1(\result[5]_i_4_n_0 ),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(memory_reg_0_i_2_n_0),
        .I5(literal_2[5]),
        .O(\result[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0C000A00))
    \result[5]_i_4
       (.I0(DATA[5]),
        .I1(OUT1[5]),
        .I2(\state_reg_n_0_[0] ),
        .I3(\state_reg_n_0_[1] ),
        .I4(read_input[1]),
        .O(\result[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[6]_i_1
       (.I0(\result[6]_i_2_n_0 ),
        .I1(\result_reg[7]_i_3_n_5 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result[6]_i_3_n_0 ),
        .I4(\result[7]_i_5_n_0 ),
        .I5(data5[6]),
        .O(\result[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00F0444400004444))
    \result[6]_i_2
       (.I0(\state_reg_n_0_[1] ),
        .I1(load_data[6]),
        .I2(data4[6]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[3]),
        .O(\result[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEECFCCCCEECCCCCC))
    \result[6]_i_3
       (.I0(data2[6]),
        .I1(\result[6]_i_4_n_0 ),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(memory_reg_0_i_2_n_0),
        .I5(literal_2[6]),
        .O(\result[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0C000A00))
    \result[6]_i_4
       (.I0(DATA[6]),
        .I1(OUT1[6]),
        .I2(\state_reg_n_0_[0] ),
        .I3(\state_reg_n_0_[1] ),
        .I4(read_input[1]),
        .O(\result[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA))
    \result[7]_i_1
       (.I0(\result[7]_i_2_n_0 ),
        .I1(\result_reg[7]_i_3_n_4 ),
        .I2(\result[16]_i_3_n_0 ),
        .I3(\result[7]_i_4_n_0 ),
        .I4(\result[7]_i_5_n_0 ),
        .I5(data5[7]),
        .O(\result[7]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[7]_i_10
       (.I0(register_a[4]),
        .I1(operand_a1),
        .I2(result[4]),
        .I3(literal_2[4]),
        .O(\result[7]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h0C000A00))
    \result[7]_i_11
       (.I0(DATA[7]),
        .I1(OUT1[7]),
        .I2(\state_reg_n_0_[0] ),
        .I3(\state_reg_n_0_[1] ),
        .I4(read_input[1]),
        .O(\result[7]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[7]_i_12
       (.I0(register_a[7]),
        .I1(operand_a1),
        .I2(register_b[7]),
        .I3(operand_b1),
        .I4(result[7]),
        .O(\result[7]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[7]_i_13
       (.I0(register_a[6]),
        .I1(operand_a1),
        .I2(register_b[6]),
        .I3(operand_b1),
        .I4(result[6]),
        .O(\result[7]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[7]_i_14
       (.I0(register_a[5]),
        .I1(operand_a1),
        .I2(register_b[5]),
        .I3(operand_b1),
        .I4(result[5]),
        .O(\result[7]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h111E22D2))
    \result[7]_i_15
       (.I0(register_a[4]),
        .I1(operand_a1),
        .I2(register_b[4]),
        .I3(operand_b1),
        .I4(result[4]),
        .O(\result[7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00F0444400004444))
    \result[7]_i_2
       (.I0(\state_reg_n_0_[1] ),
        .I1(load_data[7]),
        .I2(data4[7]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[0] ),
        .I5(opcode_2[3]),
        .O(\result[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEECFCCCCEECCCCCC))
    \result[7]_i_4
       (.I0(data2[7]),
        .I1(\result[7]_i_11_n_0 ),
        .I2(opcode_2[0]),
        .I3(opcode_2[1]),
        .I4(memory_reg_0_i_2_n_0),
        .I5(literal_2[7]),
        .O(\result[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h80))
    \result[7]_i_5
       (.I0(opcode_2[3]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[2]),
        .O(\result[7]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[7]_i_7
       (.I0(register_a[7]),
        .I1(operand_a1),
        .I2(result[7]),
        .I3(literal_2[7]),
        .O(\result[7]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[7]_i_8
       (.I0(register_a[6]),
        .I1(operand_a1),
        .I2(result[6]),
        .I3(literal_2[6]),
        .O(\result[7]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h1DE2))
    \result[7]_i_9
       (.I0(register_a[5]),
        .I1(operand_a1),
        .I2(result[5]),
        .I3(literal_2[5]),
        .O(\result[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF8000))
    \result[8]_i_1
       (.I0(opcode_2[2]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[3]),
        .I3(data5[8]),
        .I4(\result[8]_i_2_n_0 ),
        .I5(\result[8]_i_3_n_0 ),
        .O(\result[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000AC000000A000))
    \result[8]_i_2
       (.I0(data4[8]),
        .I1(data2[8]),
        .I2(opcode_2[3]),
        .I3(\state_reg_n_0_[0] ),
        .I4(opcode_2[2]),
        .I5(opcode_2[1]),
        .O(\result[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF222F222F222))
    \result[8]_i_3
       (.I0(load_data[8]),
        .I1(\result[11]_i_3_n_0 ),
        .I2(\result[9]_i_9_n_0 ),
        .I3(literal_2[8]),
        .I4(\result_reg[11]_i_5_n_7 ),
        .I5(\result[16]_i_3_n_0 ),
        .O(\result[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF8000))
    \result[9]_i_1
       (.I0(opcode_2[2]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[3]),
        .I3(data5[9]),
        .I4(\result[9]_i_3_n_0 ),
        .I5(\result[9]_i_4_n_0 ),
        .O(\result[9]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000AC000000A000))
    \result[9]_i_3
       (.I0(data4[9]),
        .I1(data2[9]),
        .I2(opcode_2[3]),
        .I3(\state_reg_n_0_[0] ),
        .I4(opcode_2[2]),
        .I5(opcode_2[1]),
        .O(\result[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF222F222F222))
    \result[9]_i_4
       (.I0(load_data[9]),
        .I1(\result[11]_i_3_n_0 ),
        .I2(\result[9]_i_9_n_0 ),
        .I3(literal_2[9]),
        .I4(\result_reg[11]_i_5_n_6 ),
        .I5(\result[16]_i_3_n_0 ),
        .O(\result[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[9]_i_5
       (.I0(result[11]),
        .I1(operand_b1),
        .I2(register_b[11]),
        .I3(operand_a1),
        .I4(register_a[11]),
        .O(\result[9]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[9]_i_6
       (.I0(result[10]),
        .I1(operand_b1),
        .I2(register_b[10]),
        .I3(operand_a1),
        .I4(register_a[10]),
        .O(\result[9]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[9]_i_7
       (.I0(result[9]),
        .I1(operand_b1),
        .I2(register_b[9]),
        .I3(operand_a1),
        .I4(register_a[9]),
        .O(\result[9]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h124712B8))
    \result[9]_i_8
       (.I0(result[8]),
        .I1(operand_b1),
        .I2(register_b[8]),
        .I3(operand_a1),
        .I4(register_a[8]),
        .O(\result[9]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00000004))
    \result[9]_i_9
       (.I0(opcode_2[3]),
        .I1(\state_reg_n_0_[0] ),
        .I2(opcode_2[2]),
        .I3(opcode_2[1]),
        .I4(opcode_2[0]),
        .O(\result[9]_i_9_n_0 ));
  FDRE \result_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[0]_i_1_n_0 ),
        .Q(result[0]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[0]_i_11
       (.CI(1'b0),
        .CO({\result_reg[0]_i_11_n_0 ,\NLW_result_reg[0]_i_11_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b1),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(\NLW_result_reg[0]_i_11_O_UNCONNECTED [3:0]),
        .S({\result[0]_i_16_n_0 ,\result[0]_i_17_n_0 ,\result[0]_i_18_n_0 ,\result[0]_i_19_n_0 }));
  CARRY4 \result_reg[0]_i_4
       (.CI(\result_reg[0]_i_7_n_0 ),
        .CO({\NLW_result_reg[0]_i_4_CO_UNCONNECTED [3],\result_reg[0]_i_4_n_1 ,\NLW_result_reg[0]_i_4_CO_UNCONNECTED [1:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(\NLW_result_reg[0]_i_4_O_UNCONNECTED [3:0]),
        .S({1'b0,\result[0]_i_8_n_0 ,\result[0]_i_9_n_0 ,\result[0]_i_10_n_0 }));
  CARRY4 \result_reg[0]_i_7
       (.CI(\result_reg[0]_i_11_n_0 ),
        .CO({\result_reg[0]_i_7_n_0 ,\NLW_result_reg[0]_i_7_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(\NLW_result_reg[0]_i_7_O_UNCONNECTED [3:0]),
        .S({\result[0]_i_12_n_0 ,\result[0]_i_13_n_0 ,\result[0]_i_14_n_0 ,\result[0]_i_15_n_0 }));
  FDRE \result_reg[10]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[10]_i_1_n_0 ),
        .Q(result[10]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[11]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[11]_i_1_n_0 ),
        .Q(result[11]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[11]_i_4
       (.CI(\result_reg[11]_i_6_n_0 ),
        .CO({\result_reg[11]_i_4_n_0 ,\NLW_result_reg[11]_i_4_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 }),
        .O(data4[11:8]),
        .S({\result[11]_i_7_n_0 ,\result[11]_i_8_n_0 ,\result[11]_i_9_n_0 ,\result[11]_i_10_n_0 }));
  CARRY4 \result_reg[11]_i_5
       (.CI(\result_reg[7]_i_3_n_0 ),
        .CO({\result_reg[11]_i_5_n_0 ,\NLW_result_reg[11]_i_5_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 }),
        .O({\result_reg[11]_i_5_n_4 ,\result_reg[11]_i_5_n_5 ,\result_reg[11]_i_5_n_6 ,\result_reg[11]_i_5_n_7 }),
        .S({\result[11]_i_11_n_0 ,\result[11]_i_12_n_0 ,\result[11]_i_13_n_0 ,\result[11]_i_14_n_0 }));
  CARRY4 \result_reg[11]_i_6
       (.CI(\result_reg[3]_i_6_n_0 ),
        .CO({\result_reg[11]_i_6_n_0 ,\NLW_result_reg[11]_i_6_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 }),
        .O(data4[7:4]),
        .S({\result[11]_i_15_n_0 ,\result[11]_i_16_n_0 ,\result[11]_i_17_n_0 ,\result[11]_i_18_n_0 }));
  FDRE \result_reg[12]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[12]_i_1_n_0 ),
        .Q(result[12]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[12]_i_3
       (.CI(\result_reg[8]_i_4_n_0 ),
        .CO({\result_reg[12]_i_3_n_0 ,\NLW_result_reg[12]_i_3_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(data2[12:9]),
        .S(program_counter_2[12:9]));
  FDRE \result_reg[13]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[13]_i_1_n_0 ),
        .Q(result[13]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[14]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[14]_i_1_n_0 ),
        .Q(result[14]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[15]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[15]_i_1_n_0 ),
        .Q(result[15]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[15]_i_2
       (.CI(\result_reg[11]_i_4_n_0 ),
        .CO({\result_reg[15]_i_2_n_0 ,\NLW_result_reg[15]_i_2_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[15]_i_1_n_0 ,\write_output[14]_i_1_n_0 ,\write_output[13]_i_1_n_0 ,\write_output[12]_i_1_n_0 }),
        .O(data4[15:12]),
        .S({\result[15]_i_4_n_0 ,\result[15]_i_5_n_0 ,\result[15]_i_6_n_0 ,\result[15]_i_7_n_0 }));
  FDRE \result_reg[16]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[16]_i_1_n_0 ),
        .Q(result[16]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[16]_i_4
       (.CI(\result_reg[16]_i_9_n_0 ),
        .CO({\result_reg[16]_i_4_n_0 ,\NLW_result_reg[16]_i_4_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O({\result_reg[16]_i_4_n_4 ,\result_reg[16]_i_4_n_5 ,\result_reg[16]_i_4_n_6 ,\result_reg[16]_i_4_n_7 }),
        .S({\result[16]_i_10_n_0 ,\result[16]_i_11_n_0 ,\result[16]_i_12_n_0 ,\result[16]_i_13_n_0 }));
  CARRY4 \result_reg[16]_i_6
       (.CI(\result_reg[15]_i_2_n_0 ),
        .CO({\result_reg[16]_i_6_n_0 ,\NLW_result_reg[16]_i_6_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[19]_i_1_n_0 ,\write_output[18]_i_1_n_0 ,\write_output[17]_i_1_n_0 ,\write_output[16]_i_1_n_0 }),
        .O(data4[19:16]),
        .S({\result[16]_i_14_n_0 ,\result[16]_i_15_n_0 ,\result[16]_i_16_n_0 ,\result[16]_i_17_n_0 }));
  CARRY4 \result_reg[16]_i_8
       (.CI(\result_reg[12]_i_3_n_0 ),
        .CO({data2[16],\NLW_result_reg[16]_i_8_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O({\NLW_result_reg[16]_i_8_O_UNCONNECTED [3],data2[15:13]}),
        .S({1'b1,program_counter_2[15:13]}));
  CARRY4 \result_reg[16]_i_9
       (.CI(\result_reg[11]_i_5_n_0 ),
        .CO({\result_reg[16]_i_9_n_0 ,\NLW_result_reg[16]_i_9_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[15]_i_1_n_0 ,\write_output[14]_i_1_n_0 ,\write_output[13]_i_1_n_0 ,\write_output[12]_i_1_n_0 }),
        .O({\result_reg[16]_i_9_n_4 ,\result_reg[16]_i_9_n_5 ,\result_reg[16]_i_9_n_6 ,\result_reg[16]_i_9_n_7 }),
        .S({\result[16]_i_21_n_0 ,\result[16]_i_22_n_0 ,\result[16]_i_23_n_0 ,\result[16]_i_24_n_0 }));
  FDRE \result_reg[17]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[17]_i_1_n_0 ),
        .Q(result[17]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[18]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[18]_i_1_n_0 ),
        .Q(result[18]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[19]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[19]_i_1_n_0 ),
        .Q(result[19]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[19]_i_2
       (.CI(\result_reg[19]_i_4_n_0 ),
        .CO({\result_reg[19]_i_2_n_0 ,\NLW_result_reg[19]_i_2_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[19]_i_1_n_0 ,\write_output[18]_i_1_n_0 ,\write_output[17]_i_1_n_0 ,\write_output[16]_i_1_n_0 }),
        .O(data5[19:16]),
        .S({\result[19]_i_5_n_0 ,\result[19]_i_6_n_0 ,\result[19]_i_7_n_0 ,\result[19]_i_8_n_0 }));
  CARRY4 \result_reg[19]_i_4
       (.CI(\result_reg[9]_i_2_n_0 ),
        .CO({\result_reg[19]_i_4_n_0 ,\NLW_result_reg[19]_i_4_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[15]_i_1_n_0 ,\write_output[14]_i_1_n_0 ,\write_output[13]_i_1_n_0 ,\write_output[12]_i_1_n_0 }),
        .O(data5[15:12]),
        .S({\result[19]_i_9_n_0 ,\result[19]_i_10_n_0 ,\result[19]_i_11_n_0 ,\result[19]_i_12_n_0 }));
  FDRE \result_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[1]_i_1_n_0 ),
        .Q(result[1]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[20]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[20]_i_1_n_0 ),
        .Q(result[20]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[21]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[21]_i_1_n_0 ),
        .Q(result[21]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[22]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[22]_i_1_n_0 ),
        .Q(result[22]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[23]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[23]_i_1_n_0 ),
        .Q(result[23]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[23]_i_2
       (.CI(\result_reg[19]_i_2_n_0 ),
        .CO({\result_reg[23]_i_2_n_0 ,\NLW_result_reg[23]_i_2_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[23]_i_1_n_0 ,\write_output[22]_i_1_n_0 ,\write_output[21]_i_1_n_0 ,\write_output[20]_i_1_n_0 }),
        .O(data5[23:20]),
        .S({\result[23]_i_4_n_0 ,\result[23]_i_5_n_0 ,\result[23]_i_6_n_0 ,\result[23]_i_7_n_0 }));
  CARRY4 \result_reg[23]_i_8
       (.CI(\result_reg[16]_i_6_n_0 ),
        .CO({\result_reg[23]_i_8_n_0 ,\NLW_result_reg[23]_i_8_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[23]_i_1_n_0 ,\write_output[22]_i_1_n_0 ,\write_output[21]_i_1_n_0 ,\write_output[20]_i_1_n_0 }),
        .O(data4[23:20]),
        .S({\result[23]_i_10_n_0 ,\result[23]_i_11_n_0 ,\result[23]_i_12_n_0 ,\result[23]_i_13_n_0 }));
  CARRY4 \result_reg[23]_i_9
       (.CI(\result_reg[16]_i_4_n_0 ),
        .CO({\result_reg[23]_i_9_n_0 ,\NLW_result_reg[23]_i_9_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O({\result_reg[23]_i_9_n_4 ,\result_reg[23]_i_9_n_5 ,\result_reg[23]_i_9_n_6 ,\result_reg[23]_i_9_n_7 }),
        .S({\result[23]_i_14_n_0 ,\result[23]_i_15_n_0 ,\result[23]_i_16_n_0 ,\result[23]_i_17_n_0 }));
  FDRE \result_reg[24]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[24]_i_1_n_0 ),
        .Q(result[24]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[25]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[25]_i_1_n_0 ),
        .Q(result[25]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[26]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[26]_i_1_n_0 ),
        .Q(result[26]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[27]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[27]_i_1_n_0 ),
        .Q(result[27]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[27]_i_2
       (.CI(\result_reg[23]_i_2_n_0 ),
        .CO({\result_reg[27]_i_2_n_0 ,\NLW_result_reg[27]_i_2_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[27]_i_1_n_0 ,\write_output[26]_i_1_n_0 ,\write_output[25]_i_1_n_0 ,\write_output[24]_i_1_n_0 }),
        .O(data5[27:24]),
        .S({\result[27]_i_4_n_0 ,\result[27]_i_5_n_0 ,\result[27]_i_6_n_0 ,\result[27]_i_7_n_0 }));
  CARRY4 \result_reg[27]_i_8
       (.CI(\result_reg[23]_i_8_n_0 ),
        .CO({\result_reg[27]_i_8_n_0 ,\NLW_result_reg[27]_i_8_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[27]_i_1_n_0 ,\write_output[26]_i_1_n_0 ,\write_output[25]_i_1_n_0 ,\write_output[24]_i_1_n_0 }),
        .O(data4[27:24]),
        .S({\result[27]_i_10_n_0 ,\result[27]_i_11_n_0 ,\result[27]_i_12_n_0 ,\result[27]_i_13_n_0 }));
  CARRY4 \result_reg[27]_i_9
       (.CI(\result_reg[23]_i_9_n_0 ),
        .CO({\result_reg[27]_i_9_n_0 ,\NLW_result_reg[27]_i_9_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O({\result_reg[27]_i_9_n_4 ,\result_reg[27]_i_9_n_5 ,\result_reg[27]_i_9_n_6 ,\result_reg[27]_i_9_n_7 }),
        .S({\result[27]_i_14_n_0 ,\result[27]_i_15_n_0 ,\result[27]_i_16_n_0 ,\result[27]_i_17_n_0 }));
  FDRE \result_reg[28]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[28]_i_1_n_0 ),
        .Q(result[28]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[29]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[29]_i_1_n_0 ),
        .Q(result[29]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[2]_i_1_n_0 ),
        .Q(result[2]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[30]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[30]_i_1_n_0 ),
        .Q(result[30]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[31]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[31]_i_2_n_0 ),
        .Q(result[31]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[31]_i_16
       (.CI(\result_reg[27]_i_8_n_0 ),
        .CO(\NLW_result_reg[31]_i_16_CO_UNCONNECTED [3:0]),
        .CYINIT(1'b0),
        .DI({1'b0,\write_output[30]_i_1_n_0 ,\write_output[29]_i_1_n_0 ,\write_output[28]_i_1_n_0 }),
        .O(data4[31:28]),
        .S({\result[31]_i_24_n_0 ,\result[31]_i_25_n_0 ,\result[31]_i_26_n_0 ,\result[31]_i_27_n_0 }));
  CARRY4 \result_reg[31]_i_17
       (.CI(\result_reg[27]_i_9_n_0 ),
        .CO(\NLW_result_reg[31]_i_17_CO_UNCONNECTED [3:0]),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O({\result_reg[31]_i_17_n_4 ,\result_reg[31]_i_17_n_5 ,\result_reg[31]_i_17_n_6 ,\result_reg[31]_i_17_n_7 }),
        .S({\result[31]_i_28_n_0 ,\result[31]_i_29_n_0 ,\result[31]_i_30_n_0 ,\result[31]_i_31_n_0 }));
  CARRY4 \result_reg[31]_i_8
       (.CI(\result_reg[27]_i_2_n_0 ),
        .CO(\NLW_result_reg[31]_i_8_CO_UNCONNECTED [3:0]),
        .CYINIT(1'b0),
        .DI({1'b0,\write_output[30]_i_1_n_0 ,\write_output[29]_i_1_n_0 ,\write_output[28]_i_1_n_0 }),
        .O(data5[31:28]),
        .S({\result[31]_i_12_n_0 ,\result[31]_i_13_n_0 ,\result[31]_i_14_n_0 ,\result[31]_i_15_n_0 }));
  FDRE \result_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[3]_i_1_n_0 ),
        .Q(result[3]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[3]_i_3
       (.CI(1'b0),
        .CO({\result_reg[3]_i_3_n_0 ,\NLW_result_reg[3]_i_3_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 }),
        .O({\result_reg[3]_i_3_n_4 ,\result_reg[3]_i_3_n_5 ,\result_reg[3]_i_3_n_6 ,\result_reg[3]_i_3_n_7 }),
        .S({\result[3]_i_7_n_0 ,\result[3]_i_8_n_0 ,\result[3]_i_9_n_0 ,\result[3]_i_10_n_0 }));
  CARRY4 \result_reg[3]_i_5
       (.CI(1'b0),
        .CO({\result_reg[3]_i_5_n_0 ,\NLW_result_reg[3]_i_5_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 }),
        .O(data5[3:0]),
        .S({\result[3]_i_12_n_0 ,\result[3]_i_13_n_0 ,\result[3]_i_14_n_0 ,\result[3]_i_15_n_0 }));
  CARRY4 \result_reg[3]_i_6
       (.CI(1'b0),
        .CO({\result_reg[3]_i_6_n_0 ,\NLW_result_reg[3]_i_6_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b1),
        .DI({\write_output[3]_i_1_n_0 ,\write_output[2]_i_1_n_0 ,\write_output[1]_i_1_n_0 ,\write_output[0]_i_1_n_0 }),
        .O(data4[3:0]),
        .S({\result[3]_i_16_n_0 ,\result[3]_i_17_n_0 ,\result[3]_i_18_n_0 ,\result[3]_i_19_n_0 }));
  FDRE \result_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[4]_i_1_n_0 ),
        .Q(result[4]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[4]_i_4
       (.CI(1'b0),
        .CO({\result_reg[4]_i_4_n_0 ,\NLW_result_reg[4]_i_4_CO_UNCONNECTED [2:0]}),
        .CYINIT(program_counter_2[0]),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(data2[4:1]),
        .S(program_counter_2[4:1]));
  FDRE \result_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[5]_i_1_n_0 ),
        .Q(result[5]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[6]_i_1_n_0 ),
        .Q(result[6]),
        .R(INTERNAL_RST_reg));
  FDRE \result_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[7]_i_1_n_0 ),
        .Q(result[7]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[7]_i_3
       (.CI(\result_reg[3]_i_3_n_0 ),
        .CO({\result_reg[7]_i_3_n_0 ,\NLW_result_reg[7]_i_3_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 }),
        .O({\result_reg[7]_i_3_n_4 ,\result_reg[7]_i_3_n_5 ,\result_reg[7]_i_3_n_6 ,\result_reg[7]_i_3_n_7 }),
        .S({\result[7]_i_7_n_0 ,\result[7]_i_8_n_0 ,\result[7]_i_9_n_0 ,\result[7]_i_10_n_0 }));
  CARRY4 \result_reg[7]_i_6
       (.CI(\result_reg[3]_i_5_n_0 ),
        .CO({\result_reg[7]_i_6_n_0 ,\NLW_result_reg[7]_i_6_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[7]_i_1_n_0 ,\write_output[6]_i_1_n_0 ,\write_output[5]_i_1_n_0 ,\write_output[4]_i_1_n_0 }),
        .O(data5[7:4]),
        .S({\result[7]_i_12_n_0 ,\result[7]_i_13_n_0 ,\result[7]_i_14_n_0 ,\result[7]_i_15_n_0 }));
  FDRE \result_reg[8]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[8]_i_1_n_0 ),
        .Q(result[8]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[8]_i_4
       (.CI(\result_reg[4]_i_4_n_0 ),
        .CO({\result_reg[8]_i_4_n_0 ,\NLW_result_reg[8]_i_4_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({1'b0,1'b0,1'b0,1'b0}),
        .O(data2[8:5]),
        .S(program_counter_2[8:5]));
  FDRE \result_reg[9]
       (.C(ETH_CLK_OBUF),
        .CE(\result[31]_i_1_n_0 ),
        .D(\result[9]_i_1_n_0 ),
        .Q(result[9]),
        .R(INTERNAL_RST_reg));
  CARRY4 \result_reg[9]_i_2
       (.CI(\result_reg[7]_i_6_n_0 ),
        .CO({\result_reg[9]_i_2_n_0 ,\NLW_result_reg[9]_i_2_CO_UNCONNECTED [2:0]}),
        .CYINIT(1'b0),
        .DI({\write_output[11]_i_1_n_0 ,\write_output[10]_i_1_n_0 ,\write_output[9]_i_1_n_0 ,\write_output[8]_i_1_n_0 }),
        .O(data5[11:8]),
        .S({\result[9]_i_5_n_0 ,\result[9]_i_6_n_0 ,\result[9]_i_7_n_0 ,\result[9]_i_8_n_0 }));
  LUT6 #(
    .INIT(64'hFFFFF7FF00000C00))
    \s_input_ps2_ack[0]_i_1
       (.I0(S_DATA_STB_reg_0),
        .I1(\result[31]_i_3_n_0 ),
        .I2(read_input[1]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\state_reg_n_0_[0] ),
        .I5(DATA_ACK),
        .O(\s_input_ps2_ack[0]_i_1_n_0 ));
  FDRE \s_input_ps2_ack_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(1'b1),
        .D(\s_input_ps2_ack[0]_i_1_n_0 ),
        .Q(DATA_ACK),
        .R(INTERNAL_RST_reg));
  LUT6 #(
    .INIT(64'hFFFF7FFF0000C000))
    \s_input_rs232_rx_ack[0]_i_1
       (.I0(OUT1_STB),
        .I1(\result[31]_i_3_n_0 ),
        .I2(read_input[1]),
        .I3(\state_reg_n_0_[1] ),
        .I4(\state_reg_n_0_[0] ),
        .I5(OUT1_ACK),
        .O(\s_input_rs232_rx_ack[0]_i_1_n_0 ));
  FDRE \s_input_rs232_rx_ack_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(1'b1),
        .D(\s_input_rs232_rx_ack[0]_i_1_n_0 ),
        .Q(OUT1_ACK),
        .R(INTERNAL_RST_reg));
  LUT6 #(
    .INIT(64'h0000000200000000))
    \s_output_rs232_tx[7]_i_1
       (.I0(\s_output_rs232_tx[7]_i_2_n_0 ),
        .I1(write_output[13]),
        .I2(write_output[12]),
        .I3(write_output[15]),
        .I4(write_output[14]),
        .I5(\s_output_rs232_tx[7]_i_3_n_0 ),
        .O(E));
  LUT6 #(
    .INIT(64'h0000000000008000))
    \s_output_rs232_tx[7]_i_2
       (.I0(\s_output_rs232_tx[7]_i_4_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(\state_reg_n_0_[1] ),
        .I3(\state_reg_n_0_[2] ),
        .I4(write_output[8]),
        .I5(write_output[9]),
        .O(\s_output_rs232_tx[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000002000000000))
    \s_output_rs232_tx[7]_i_3
       (.I0(\s_output_rs232_tx[7]_i_5_n_0 ),
        .I1(write_output[1]),
        .I2(write_output[0]),
        .I3(write_output[3]),
        .I4(write_output[2]),
        .I5(\s_output_rs232_tx[7]_i_6_n_0 ),
        .O(\s_output_rs232_tx[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0001))
    \s_output_rs232_tx[7]_i_4
       (.I0(write_output[5]),
        .I1(write_output[4]),
        .I2(write_output[7]),
        .I3(write_output[6]),
        .O(\s_output_rs232_tx[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001))
    \s_output_rs232_tx[7]_i_5
       (.I0(write_output[29]),
        .I1(write_output[28]),
        .I2(write_output[22]),
        .I3(write_output[23]),
        .I4(write_output[30]),
        .I5(write_output[31]),
        .O(\s_output_rs232_tx[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8))
    \s_output_rs232_tx[7]_i_6
       (.I0(\s_output_rs232_tx[7]_i_7_n_0 ),
        .I1(\s_output_rs232_tx[7]_i_8_n_0 ),
        .O(\s_output_rs232_tx[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001))
    \s_output_rs232_tx[7]_i_7
       (.I0(write_output[19]),
        .I1(write_output[18]),
        .I2(write_output[10]),
        .I3(write_output[11]),
        .I4(write_output[20]),
        .I5(write_output[21]),
        .O(\s_output_rs232_tx[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001))
    \s_output_rs232_tx[7]_i_8
       (.I0(write_output[25]),
        .I1(write_output[24]),
        .I2(write_output[16]),
        .I3(write_output[17]),
        .I4(write_output[26]),
        .I5(write_output[27]),
        .O(\s_output_rs232_tx[7]_i_8_n_0 ));
  FDRE \s_output_rs232_tx_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(E),
        .D(write_value[0]),
        .Q(Q[0]),
        .R(1'b0));
  FDRE \s_output_rs232_tx_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(E),
        .D(write_value[1]),
        .Q(Q[1]),
        .R(1'b0));
  FDRE \s_output_rs232_tx_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(E),
        .D(write_value[2]),
        .Q(Q[2]),
        .R(1'b0));
  FDRE \s_output_rs232_tx_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(E),
        .D(write_value[3]),
        .Q(Q[3]),
        .R(1'b0));
  FDRE \s_output_rs232_tx_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(E),
        .D(write_value[4]),
        .Q(Q[4]),
        .R(1'b0));
  FDRE \s_output_rs232_tx_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(E),
        .D(write_value[5]),
        .Q(Q[5]),
        .R(1'b0));
  FDRE \s_output_rs232_tx_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(E),
        .D(write_value[6]),
        .Q(Q[6]),
        .R(1'b0));
  FDRE \s_output_rs232_tx_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(E),
        .D(write_value[7]),
        .Q(Q[7]),
        .R(1'b0));
  FDRE \s_output_rs232_tx_stb_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(1'b1),
        .D(S_IN1_ACK_reg),
        .Q(IN1_STB),
        .R(INTERNAL_RST_reg));
  LUT6 #(
    .INIT(64'hEAFAFFFFFAFA0000))
    \state[0]_i_1
       (.I0(\state_reg_n_0_[2] ),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[1] ),
        .I3(opcode_2[2]),
        .I4(\state[2]_i_3_n_0 ),
        .I5(\state_reg_n_0_[0] ),
        .O(\state[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFDDDFFFFFFFF0000))
    \state[1]_i_1
       (.I0(\state_reg_n_0_[0] ),
        .I1(\state_reg_n_0_[2] ),
        .I2(opcode_2[2]),
        .I3(opcode_2[1]),
        .I4(\state[2]_i_3_n_0 ),
        .I5(\state_reg_n_0_[1] ),
        .O(\state[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h88A8FFFF88A80000))
    \state[2]_i_1
       (.I0(\state[2]_i_2_n_0 ),
        .I1(opcode_2[1]),
        .I2(opcode_2[0]),
        .I3(opcode_2[3]),
        .I4(\state[2]_i_3_n_0 ),
        .I5(\state_reg_n_0_[2] ),
        .O(\state[2]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8000))
    \state[2]_i_10
       (.I0(\state[2]_i_13_n_0 ),
        .I1(\s_output_rs232_tx[7]_i_6_n_0 ),
        .I2(\state[2]_i_14_n_0 ),
        .I3(\state[2]_i_15_n_0 ),
        .O(\state[2]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hAFBE))
    \state[2]_i_11
       (.I0(\state[2]_i_16_n_0 ),
        .I1(\state_reg_n_0_[0] ),
        .I2(\state_reg_n_0_[1] ),
        .I3(\state_reg_n_0_[2] ),
        .O(\state[2]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h08000000))
    \state[2]_i_12
       (.I0(read_input[1]),
        .I1(\state_reg_n_0_[1] ),
        .I2(\state_reg_n_0_[0] ),
        .I3(OUT1_ACK),
        .I4(OUT1_STB),
        .O(\state[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000))
    \state[2]_i_13
       (.I0(\state[2]_i_17_n_0 ),
        .I1(write_output[9]),
        .I2(write_output[8]),
        .I3(\state_reg_n_0_[2] ),
        .I4(\state_reg_n_0_[0] ),
        .I5(\s_output_rs232_tx[7]_i_4_n_0 ),
        .O(\state[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004))
    \state[2]_i_14
       (.I0(write_output[1]),
        .I1(write_output[0]),
        .I2(write_output[28]),
        .I3(write_output[29]),
        .I4(write_output[2]),
        .I5(write_output[3]),
        .O(\state[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000))
    \state[2]_i_15
       (.I0(write_output[31]),
        .I1(write_output[30]),
        .I2(IN1_STB),
        .I3(IN1_ACK),
        .I4(write_output[22]),
        .I5(write_output[23]),
        .O(\state[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000035400000))
    \state[2]_i_16
       (.I0(opcode_2[3]),
        .I1(opcode_2[0]),
        .I2(opcode_2[1]),
        .I3(opcode_2[2]),
        .I4(\state_reg_n_0_[1] ),
        .I5(\state_reg_n_0_[2] ),
        .O(\state[2]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0001))
    \state[2]_i_17
       (.I0(write_output[13]),
        .I1(write_output[12]),
        .I2(write_output[15]),
        .I3(write_output[14]),
        .O(\state[2]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0080))
    \state[2]_i_2
       (.I0(\state_reg_n_0_[0] ),
        .I1(opcode_2[2]),
        .I2(\state_reg_n_0_[1] ),
        .I3(\state_reg_n_0_[2] ),
        .O(\state[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF30FFB0FFB0))
    \state[2]_i_3
       (.I0(\state[2]_i_4_n_0 ),
        .I1(\state[2]_i_5_n_0 ),
        .I2(\state[2]_i_6_n_0 ),
        .I3(\state[2]_i_7_n_0 ),
        .I4(\state[2]_i_8_n_0 ),
        .I5(\program_counter_rep[9]_i_7_n_0 ),
        .O(\state[2]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1))
    \state[2]_i_4
       (.I0(opcode_2[1]),
        .I1(opcode_2[2]),
        .O(\state[2]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hB))
    \state[2]_i_5
       (.I0(opcode_2[1]),
        .I1(opcode_2[0]),
        .O(\state[2]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h08))
    \state[2]_i_6
       (.I0(\state_reg_n_0_[1] ),
        .I1(opcode_2[3]),
        .I2(\state_reg_n_0_[2] ),
        .O(\state[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF4FFF0FFF0))
    \state[2]_i_7
       (.I0(S_DATA_STB_reg),
        .I1(\state[2]_i_9_n_0 ),
        .I2(\state[2]_i_10_n_0 ),
        .I3(\state[2]_i_11_n_0 ),
        .I4(\state[2]_i_12_n_0 ),
        .I5(\result[31]_i_10_n_0 ),
        .O(\state[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00000080))
    \state[2]_i_8
       (.I0(opcode_2[3]),
        .I1(\state_reg_n_0_[1] ),
        .I2(opcode_2[1]),
        .I3(opcode_2[0]),
        .I4(\state_reg_n_0_[2] ),
        .O(\state[2]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h04))
    \state[2]_i_9
       (.I0(\state_reg_n_0_[0] ),
        .I1(\state_reg_n_0_[1] ),
        .I2(read_input[1]),
        .O(\state[2]_i_9_n_0 ));
  FDSE \state_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(1'b1),
        .D(\state[0]_i_1_n_0 ),
        .Q(\state_reg_n_0_[0] ),
        .S(INTERNAL_RST_reg));
  FDRE \state_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(1'b1),
        .D(\state[1]_i_1_n_0 ),
        .Q(\state_reg_n_0_[1] ),
        .R(INTERNAL_RST_reg));
  FDRE \state_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(1'b1),
        .D(\state[2]_i_1_n_0 ),
        .Q(\state_reg_n_0_[2] ),
        .R(INTERNAL_RST_reg));
  FDRE write_enable_reg
       (.C(ETH_CLK_OBUF),
        .CE(1'b1),
        .D(\result[31]_i_1_n_0 ),
        .Q(write_enable),
        .R(1'b0));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[0]_i_1
       (.I0(result[0]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[0]),
        .O(\write_output[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[10]_i_1
       (.I0(result[10]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[10]),
        .O(\write_output[10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[11]_i_1
       (.I0(result[11]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[11]),
        .O(\write_output[11]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[12]_i_1
       (.I0(result[12]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[12]),
        .O(\write_output[12]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[13]_i_1
       (.I0(result[13]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[13]),
        .O(\write_output[13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[14]_i_1
       (.I0(result[14]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[14]),
        .O(\write_output[14]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[15]_i_1
       (.I0(result[15]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[15]),
        .O(\write_output[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[16]_i_1
       (.I0(result[16]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[16]),
        .O(\write_output[16]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[17]_i_1
       (.I0(result[17]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[17]),
        .O(\write_output[17]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[18]_i_1
       (.I0(result[18]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[18]),
        .O(\write_output[18]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[19]_i_1
       (.I0(result[19]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[19]),
        .O(\write_output[19]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[1]_i_1
       (.I0(result[1]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[1]),
        .O(\write_output[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[20]_i_1
       (.I0(result[20]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[20]),
        .O(\write_output[20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[21]_i_1
       (.I0(result[21]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[21]),
        .O(\write_output[21]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[22]_i_1
       (.I0(result[22]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[22]),
        .O(\write_output[22]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[23]_i_1
       (.I0(result[23]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[23]),
        .O(\write_output[23]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[24]_i_1
       (.I0(result[24]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[24]),
        .O(\write_output[24]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[25]_i_1
       (.I0(result[25]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[25]),
        .O(\write_output[25]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[26]_i_1
       (.I0(result[26]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[26]),
        .O(\write_output[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[27]_i_1
       (.I0(result[27]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[27]),
        .O(\write_output[27]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[28]_i_1
       (.I0(result[28]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[28]),
        .O(\write_output[28]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[29]_i_1
       (.I0(result[29]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[29]),
        .O(\write_output[29]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[2]_i_1
       (.I0(result[2]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[2]),
        .O(\write_output[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[30]_i_1
       (.I0(result[30]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[30]),
        .O(\write_output[30]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000000))
    \write_output[31]_i_1
       (.I0(\state_reg_n_0_[2] ),
        .I1(\write_output[31]_i_3_n_0 ),
        .I2(opcode_2[3]),
        .I3(\state_reg_n_0_[1] ),
        .I4(opcode_2[1]),
        .I5(opcode_2[0]),
        .O(\write_output[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[31]_i_2
       (.I0(result[31]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[31]),
        .O(\write_output[31]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7))
    \write_output[31]_i_3
       (.I0(opcode_2[2]),
        .I1(\state_reg_n_0_[0] ),
        .O(\write_output[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009))
    \write_output[31]_i_4
       (.I0(address_a_2[2]),
        .I1(address_z_3[2]),
        .I2(address_a_2[1]),
        .I3(address_z_3[1]),
        .I4(address_z_3[0]),
        .I5(address_a_2[0]),
        .O(\write_output[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[3]_i_1
       (.I0(result[3]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[3]),
        .O(\write_output[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[4]_i_1
       (.I0(result[4]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[4]),
        .O(\write_output[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[5]_i_1
       (.I0(result[5]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[5]),
        .O(\write_output[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[6]_i_1
       (.I0(result[6]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[6]),
        .O(\write_output[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[7]_i_1
       (.I0(result[7]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[7]),
        .O(\write_output[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[8]_i_1
       (.I0(result[8]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[8]),
        .O(\write_output[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFBF80000080))
    \write_output[9]_i_1
       (.I0(result[9]),
        .I1(\write_output[31]_i_4_n_0 ),
        .I2(write_enable),
        .I3(address_a_2[3]),
        .I4(address_z_3[3]),
        .I5(register_a[9]),
        .O(\write_output[9]_i_1_n_0 ));
  FDRE \write_output_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[0]_i_1_n_0 ),
        .Q(write_output[0]),
        .R(1'b0));
  FDRE \write_output_reg[10]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[10]_i_1_n_0 ),
        .Q(write_output[10]),
        .R(1'b0));
  FDRE \write_output_reg[11]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[11]_i_1_n_0 ),
        .Q(write_output[11]),
        .R(1'b0));
  FDRE \write_output_reg[12]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[12]_i_1_n_0 ),
        .Q(write_output[12]),
        .R(1'b0));
  FDRE \write_output_reg[13]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[13]_i_1_n_0 ),
        .Q(write_output[13]),
        .R(1'b0));
  FDRE \write_output_reg[14]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[14]_i_1_n_0 ),
        .Q(write_output[14]),
        .R(1'b0));
  FDRE \write_output_reg[15]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[15]_i_1_n_0 ),
        .Q(write_output[15]),
        .R(1'b0));
  FDRE \write_output_reg[16]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[16]_i_1_n_0 ),
        .Q(write_output[16]),
        .R(1'b0));
  FDRE \write_output_reg[17]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[17]_i_1_n_0 ),
        .Q(write_output[17]),
        .R(1'b0));
  FDRE \write_output_reg[18]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[18]_i_1_n_0 ),
        .Q(write_output[18]),
        .R(1'b0));
  FDRE \write_output_reg[19]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[19]_i_1_n_0 ),
        .Q(write_output[19]),
        .R(1'b0));
  FDRE \write_output_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[1]_i_1_n_0 ),
        .Q(write_output[1]),
        .R(1'b0));
  FDRE \write_output_reg[20]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[20]_i_1_n_0 ),
        .Q(write_output[20]),
        .R(1'b0));
  FDRE \write_output_reg[21]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[21]_i_1_n_0 ),
        .Q(write_output[21]),
        .R(1'b0));
  FDRE \write_output_reg[22]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[22]_i_1_n_0 ),
        .Q(write_output[22]),
        .R(1'b0));
  FDRE \write_output_reg[23]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[23]_i_1_n_0 ),
        .Q(write_output[23]),
        .R(1'b0));
  FDRE \write_output_reg[24]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[24]_i_1_n_0 ),
        .Q(write_output[24]),
        .R(1'b0));
  FDRE \write_output_reg[25]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[25]_i_1_n_0 ),
        .Q(write_output[25]),
        .R(1'b0));
  FDRE \write_output_reg[26]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[26]_i_1_n_0 ),
        .Q(write_output[26]),
        .R(1'b0));
  FDRE \write_output_reg[27]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[27]_i_1_n_0 ),
        .Q(write_output[27]),
        .R(1'b0));
  FDRE \write_output_reg[28]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[28]_i_1_n_0 ),
        .Q(write_output[28]),
        .R(1'b0));
  FDRE \write_output_reg[29]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[29]_i_1_n_0 ),
        .Q(write_output[29]),
        .R(1'b0));
  FDRE \write_output_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[2]_i_1_n_0 ),
        .Q(write_output[2]),
        .R(1'b0));
  FDRE \write_output_reg[30]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[30]_i_1_n_0 ),
        .Q(write_output[30]),
        .R(1'b0));
  FDRE \write_output_reg[31]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[31]_i_2_n_0 ),
        .Q(write_output[31]),
        .R(1'b0));
  FDRE \write_output_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[3]_i_1_n_0 ),
        .Q(write_output[3]),
        .R(1'b0));
  FDRE \write_output_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[4]_i_1_n_0 ),
        .Q(write_output[4]),
        .R(1'b0));
  FDRE \write_output_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[5]_i_1_n_0 ),
        .Q(write_output[5]),
        .R(1'b0));
  FDRE \write_output_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[6]_i_1_n_0 ),
        .Q(write_output[6]),
        .R(1'b0));
  FDRE \write_output_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[7]_i_1_n_0 ),
        .Q(write_output[7]),
        .R(1'b0));
  FDRE \write_output_reg[8]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[8]_i_1_n_0 ),
        .Q(write_output[8]),
        .R(1'b0));
  FDRE \write_output_reg[9]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(\write_output[9]_i_1_n_0 ),
        .Q(write_output[9]),
        .R(1'b0));
  LUT3 #(
    .INIT(8'hB8))
    \write_value[0]_i_1
       (.I0(result[0]),
        .I1(operand_b1),
        .I2(register_b[0]),
        .O(store_data[0]));
  LUT3 #(
    .INIT(8'hB8))
    \write_value[1]_i_1
       (.I0(result[1]),
        .I1(operand_b1),
        .I2(register_b[1]),
        .O(store_data[1]));
  LUT3 #(
    .INIT(8'hB8))
    \write_value[2]_i_1
       (.I0(result[2]),
        .I1(operand_b1),
        .I2(register_b[2]),
        .O(store_data[2]));
  LUT3 #(
    .INIT(8'hB8))
    \write_value[3]_i_1
       (.I0(result[3]),
        .I1(operand_b1),
        .I2(register_b[3]),
        .O(store_data[3]));
  LUT3 #(
    .INIT(8'hB8))
    \write_value[4]_i_1
       (.I0(result[4]),
        .I1(operand_b1),
        .I2(register_b[4]),
        .O(store_data[4]));
  LUT3 #(
    .INIT(8'hB8))
    \write_value[5]_i_1
       (.I0(result[5]),
        .I1(operand_b1),
        .I2(register_b[5]),
        .O(store_data[5]));
  LUT3 #(
    .INIT(8'hB8))
    \write_value[6]_i_1
       (.I0(result[6]),
        .I1(operand_b1),
        .I2(register_b[6]),
        .O(store_data[6]));
  LUT3 #(
    .INIT(8'hB8))
    \write_value[7]_i_1
       (.I0(result[7]),
        .I1(operand_b1),
        .I2(register_b[7]),
        .O(store_data[7]));
  LUT4 #(
    .INIT(16'h8008))
    \write_value[7]_i_2
       (.I0(\write_value[7]_i_3_n_0 ),
        .I1(write_enable),
        .I2(address_z_3[3]),
        .I3(address_b_2[3]),
        .O(operand_b1));
  LUT6 #(
    .INIT(64'h9009000000009009))
    \write_value[7]_i_3
       (.I0(address_z_3[2]),
        .I1(address_b_2[2]),
        .I2(address_z_3[1]),
        .I3(address_b_2[1]),
        .I4(address_b_2[0]),
        .I5(address_z_3[0]),
        .O(\write_value[7]_i_3_n_0 ));
  FDRE \write_value_reg[0]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(store_data[0]),
        .Q(write_value[0]),
        .R(1'b0));
  FDRE \write_value_reg[1]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(store_data[1]),
        .Q(write_value[1]),
        .R(1'b0));
  FDRE \write_value_reg[2]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(store_data[2]),
        .Q(write_value[2]),
        .R(1'b0));
  FDRE \write_value_reg[3]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(store_data[3]),
        .Q(write_value[3]),
        .R(1'b0));
  FDRE \write_value_reg[4]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(store_data[4]),
        .Q(write_value[4]),
        .R(1'b0));
  FDRE \write_value_reg[5]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(store_data[5]),
        .Q(write_value[5]),
        .R(1'b0));
  FDRE \write_value_reg[6]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(store_data[6]),
        .Q(write_value[6]),
        .R(1'b0));
  FDRE \write_value_reg[7]
       (.C(ETH_CLK_OBUF),
        .CE(\write_output[31]_i_1_n_0 ),
        .D(store_data[7]),
        .Q(write_value[7]),
        .R(1'b0));
endmodule