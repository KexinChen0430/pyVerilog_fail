module bug98(interfacex x_if);
   h inst_h(.push(x_if.pop));
endmodule