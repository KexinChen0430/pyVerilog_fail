module test_bsg
#(
  parameter width_p      = `WIDTH_P,
  parameter cycle_time_p = 20,
  parameter reset_cycles_lo_p=0,
  parameter reset_cycles_hi_p=5
);
  wire clk;
  wire reset;
  bsg_nonsynth_clock_gen #(  .cycle_time_p(cycle_time_p)
                          )  clock_gen
                          (  .o(clk)
                          );
  bsg_nonsynth_reset_gen #(  .num_clocks_p     (1)
                           , .reset_cycles_lo_p(reset_cycles_lo_p)
                           , .reset_cycles_hi_p(reset_cycles_hi_p)
                          )  reset_gen
                          (  .clk_i        (clk)
                           , .async_reset_o(reset)
                          );
  initial
  begin
    $display("\n\n\n");
    $display("===========================================================");
    $display("testing with ...");
    $display("WIDTH_P: %d\n", width_p);
  end
  logic [width_p-1:0]           test_input, test_input_n;
  logic [width_p-1:0]           count;
  logic [$clog2(width_p+1)-1:0] test_output, popcount; //popcount is expected output
  logic finish_r;
  // Gray codes are used as test inputs since pop code of gray code of every
  // next number is incremented/decremented only once.
  if(width_p > 1)
    bsg_binary_plus_one_to_gray #(  .width_p(width_p)
                                 )  binary_pone_gray
                                 (  .binary_i(width_p'(count-1))
                                  , .gray_o  (test_input_n)
                                 );
  else
    assign test_input_n = count;
  always_ff @(posedge clk)
  begin
    test_input   <= test_input_n;
    if(reset)
      begin
        count    <= 0;
        popcount <= 0;
      end
    else
      begin
        count <= count + 1;
        if(test_input_n > test_input)
          popcount <= popcount + 1;
        else if(test_input_n < test_input)
          popcount <= popcount - 1;
      end
  end
  always_ff @(posedge clk)
  begin
    /*$display("\ncount: %b, test_input: %b, test_output: %b"
             , count, test_input, test_output);*/
    if(!reset)
      assert(test_output == popcount)
        else $error("mismatch on input %b, expected output: %b, test_output:%b"
                    , test_input, popcount, test_output);
    if(&count)
      finish_r <= 1'b1;
    if(finish_r)
      begin
        $display("=============================================================\n");
        $finish;
      end
  end
  bsg_popcount #(  .width_p(width_p)
                )  DUT
                (  .i(test_input)
                 , .o(test_output)
                );
  /*logic [(3*width_p)-1:0] log;
  assign log = {  width_p'(test_output)
                , width_p'(popcount)
                , test_input};
  bsg_nonsynth_ascii_writer #(  .width_p      (width_p)
                              , .values_p     (3)
                              , .filename_p   ("output.log")
                              , .fopen_param_p("a+")
                              , .format_p     ("%x")
                             )  ascii_writer
                             (  .clk    (clk)
                              , .reset_i(reset)
                              , .valid_i(1'b1)
                              , .data_i (log)
                             );*/
endmodule