module bsg_mesh_to_ring_stitch   #(parameter `BSG_INV_PARAM(y_max_p)
                                  ,parameter `BSG_INV_PARAM(x_max_p)
                                  ,parameter `BSG_INV_PARAM(width_back_p)
                                  ,parameter `BSG_INV_PARAM(width_fwd_p)
                                  ,parameter b_lp = $clog2(x_max_p*y_max_p)
                                  ) (output  [x_max_p-1:0][y_max_p-1:0][b_lp-1:0] id_o
                                     ,output [x_max_p-1:0][y_max_p-1:0][width_back_p-1:0] back_data_in_o
                                     ,input  [x_max_p-1:0][y_max_p-1:0][width_back_p-1:0] back_data_out_i
                                     ,output [x_max_p-1:0][y_max_p-1:0][width_fwd_p-1:0]  fwd_data_in_o
                                     ,input  [x_max_p-1:0][y_max_p-1:0][width_fwd_p-1:0]  fwd_data_out_i
                                    );
if (x_max_p == 2  && y_max_p == 2 )
begin
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  0 <- 1
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 1 ][ 1 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  3 <- 0
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  3 -> 0
 assign id_o =
 {
// y =  0,  1,
  { b_lp ' (3) , b_lp ' (0)     }, // x =  0
  { b_lp ' (2) , b_lp ' (1)     } // x =  1
 };
end
if (x_max_p == 2  && y_max_p == 3 )
begin
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 1 ][ 2 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  2 -> 3
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 1 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  5 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 0 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  4 -> 5
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  4 <- 5
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  5 -> 0
 assign id_o =
 {
// y =  0,  1,  2,
  { b_lp ' (5) , b_lp ' (0) , b_lp ' (1)     }, // x =  0
  { b_lp ' (4) , b_lp ' (3) , b_lp ' (2)     } // x =  1
 };
end
if (x_max_p == 2  && y_max_p == 4 )
begin
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 1 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  7 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 0 ]; //  5 <- 6
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  6 -> 7
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  6 <- 7
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  7 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,
  { b_lp ' (7) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2)     }, // x =  0
  { b_lp ' (6) , b_lp ' (5) , b_lp ' (4) , b_lp ' (3)     } // x =  1
 };
end
if (x_max_p == 2  && y_max_p == 5 )
begin
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 1 ][ 4 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 1 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  9 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 0 ]; //  7 <- 8
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  8 -> 9
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  8 <- 9
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  9 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,
  { b_lp ' (9) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3)     }, // x =  0
  { b_lp ' (8) , b_lp ' (7) , b_lp ' (6) , b_lp ' (5) , b_lp ' (4)     } // x =  1
 };
end
if (x_max_p == 2  && y_max_p == 6 )
begin
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 1 ][ 1 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  11 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 0 ]; //  9 <- 10
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  10 <- 11
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  11 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,
  { b_lp ' (11) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4)     }, // x =  0
  { b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7) , b_lp ' (6) , b_lp ' (5)     } // x =  1
 };
end
if (x_max_p == 2  && y_max_p == 7 )
begin
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 1 ][ 6 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 1 ][ 6 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 6 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 0 ][ 6 ]; //  5 -> 6
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 1 ][ 5 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 1 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  13 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 0 ]; //  11 <- 12
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  12 -> 13
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  12 <- 13
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  13 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,
  { b_lp ' (13) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4) , b_lp ' (5)     }, // x =  0
  { b_lp ' (12) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7) , b_lp ' (6)     } // x =  1
 };
end
if (x_max_p == 2  && y_max_p == 8 )
begin
assign back_data_in_o[ 0 ][ 7 ] = back_data_out_i[ 1 ][ 7 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 1 ][ 7 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 0 ][ 7 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 7 ] = fwd_data_out_i [ 0 ][ 7 ]; //  6 -> 7
assign back_data_in_o[ 1 ][ 7 ] = back_data_out_i[ 1 ][ 6 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 1 ][ 6 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 6 ]; //  4 <- 5
assign fwd_data_in_o [ 0 ][ 7 ] = fwd_data_out_i [ 0 ][ 6 ]; //  5 -> 6
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 1 ][ 5 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  10 -> 11
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  11 <- 12
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  12 -> 13
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  12 <- 13
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 1 ][ 1 ]; //  13 -> 14
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  15 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 0 ]; //  13 <- 14
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  14 <- 15
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  15 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,  7,
  { b_lp ' (15) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4) , b_lp ' (5) , b_lp ' (6)     }, // x =  0
  { b_lp ' (14) , b_lp ' (13) , b_lp ' (12) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7)     } // x =  1
 };
end
if (x_max_p == 4  && y_max_p == 2 )
begin
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 3 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  1 <- 2
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  2 -> 3
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  0 <- 1
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  7 <- 0
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 3 ][ 0 ]; //  3 <- 4
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  4 -> 5
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  5 -> 6
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  5 <- 6
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  6 -> 7
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  6 <- 7
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  7 -> 0
 assign id_o =
 {
// y =  0,  1,
  { b_lp ' (7) , b_lp ' (0)     }, // x =  0
  { b_lp ' (6) , b_lp ' (1)     }, // x =  1
  { b_lp ' (5) , b_lp ' (2)     }, // x =  2
  { b_lp ' (4) , b_lp ' (3)     } // x =  3
 };
end
if (x_max_p == 4  && y_max_p == 3 )
begin
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  5 <- 6
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  4 <- 5
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 1 ][ 2 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  2 -> 3
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 3 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  11 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 3 ][ 0 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  8 -> 9
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  9 -> 10
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  9 <- 10
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  10 <- 11
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  11 -> 0
 assign id_o =
 {
// y =  0,  1,  2,
  { b_lp ' (11) , b_lp ' (0) , b_lp ' (1)     }, // x =  0
  { b_lp ' (10) , b_lp ' (3) , b_lp ' (2)     }, // x =  1
  { b_lp ' (9) , b_lp ' (4) , b_lp ' (5)     }, // x =  2
  { b_lp ' (8) , b_lp ' (7) , b_lp ' (6)     } // x =  3
 };
end
if (x_max_p == 4  && y_max_p == 4 )
begin
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  8 <- 9
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  9 -> 10
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  7 <- 8
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  6 <- 7
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  7 -> 8
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 3 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  15 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 3 ][ 0 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  12 -> 13
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  12 <- 13
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  13 -> 14
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  13 <- 14
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  14 <- 15
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  15 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,
  { b_lp ' (15) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2)     }, // x =  0
  { b_lp ' (14) , b_lp ' (5) , b_lp ' (4) , b_lp ' (3)     }, // x =  1
  { b_lp ' (13) , b_lp ' (6) , b_lp ' (7) , b_lp ' (8)     }, // x =  2
  { b_lp ' (12) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9)     } // x =  3
 };
end
if (x_max_p == 4  && y_max_p == 5 )
begin
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 3 ][ 4 ]; //  11 <- 12
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  12 -> 13
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  10 <- 11
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 2 ][ 4 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 1 ][ 4 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  12 <- 13
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  13 -> 14
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  9 <- 10
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  13 <- 14
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  14 <- 15
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 3 ][ 1 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  19 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 3 ][ 0 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  16 -> 17
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  16 <- 17
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  17 -> 18
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  17 <- 18
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  18 -> 19
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  18 <- 19
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  19 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,
  { b_lp ' (19) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3)     }, // x =  0
  { b_lp ' (18) , b_lp ' (7) , b_lp ' (6) , b_lp ' (5) , b_lp ' (4)     }, // x =  1
  { b_lp ' (17) , b_lp ' (8) , b_lp ' (9) , b_lp ' (10) , b_lp ' (11)     }, // x =  2
  { b_lp ' (16) , b_lp ' (15) , b_lp ' (14) , b_lp ' (13) , b_lp ' (12)     } // x =  3
 };
end
if (x_max_p == 4  && y_max_p == 6 )
begin
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 3 ][ 5 ]; //  14 <- 15
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  15 -> 16
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  13 <- 14
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  14 -> 15
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  15 <- 16
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  16 -> 17
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  16 <- 17
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  17 -> 18
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  12 -> 13
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  17 <- 18
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  18 -> 19
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  10 <- 11
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  11 -> 12
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  18 <- 19
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 3 ][ 1 ]; //  19 -> 20
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  9 <- 10
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  23 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 3 ][ 0 ]; //  19 <- 20
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  20 -> 21
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  20 <- 21
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  21 <- 22
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  22 -> 23
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  22 <- 23
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  23 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,
  { b_lp ' (23) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4)     }, // x =  0
  { b_lp ' (22) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7) , b_lp ' (6) , b_lp ' (5)     }, // x =  1
  { b_lp ' (21) , b_lp ' (10) , b_lp ' (11) , b_lp ' (12) , b_lp ' (13) , b_lp ' (14)     }, // x =  2
  { b_lp ' (20) , b_lp ' (19) , b_lp ' (18) , b_lp ' (17) , b_lp ' (16) , b_lp ' (15)     } // x =  3
 };
end
if (x_max_p == 4  && y_max_p == 7 )
begin
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 3 ][ 6 ]; //  17 <- 18
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 3 ][ 6 ]; //  18 -> 19
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 2 ][ 6 ]; //  16 <- 17
assign fwd_data_in_o [ 3 ][ 6 ] = fwd_data_out_i [ 2 ][ 6 ]; //  17 -> 18
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 1 ][ 6 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 1 ][ 6 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 6 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 0 ][ 6 ]; //  5 -> 6
assign back_data_in_o[ 3 ][ 6 ] = back_data_out_i[ 3 ][ 5 ]; //  18 <- 19
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  19 -> 20
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 2 ][ 5 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 1 ][ 5 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  20 -> 21
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  14 <- 15
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  21 <- 22
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  22 <- 23
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 3 ][ 1 ]; //  23 -> 24
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  12 -> 13
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  27 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 3 ][ 0 ]; //  23 <- 24
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  24 -> 25
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  24 <- 25
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  25 -> 26
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  25 <- 26
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  26 -> 27
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  26 <- 27
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  27 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,
  { b_lp ' (27) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4) , b_lp ' (5)     }, // x =  0
  { b_lp ' (26) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7) , b_lp ' (6)     }, // x =  1
  { b_lp ' (25) , b_lp ' (12) , b_lp ' (13) , b_lp ' (14) , b_lp ' (15) , b_lp ' (16) , b_lp ' (17)     }, // x =  2
  { b_lp ' (24) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21) , b_lp ' (20) , b_lp ' (19) , b_lp ' (18)     } // x =  3
 };
end
if (x_max_p == 4  && y_max_p == 8 )
begin
assign back_data_in_o[ 2 ][ 7 ] = back_data_out_i[ 3 ][ 7 ]; //  20 <- 21
assign fwd_data_in_o [ 3 ][ 6 ] = fwd_data_out_i [ 3 ][ 7 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 2 ][ 7 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 7 ] = fwd_data_out_i [ 2 ][ 7 ]; //  20 -> 21
assign back_data_in_o[ 0 ][ 7 ] = back_data_out_i[ 1 ][ 7 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 1 ][ 7 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 0 ][ 7 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 7 ] = fwd_data_out_i [ 0 ][ 7 ]; //  6 -> 7
assign back_data_in_o[ 3 ][ 7 ] = back_data_out_i[ 3 ][ 6 ]; //  21 <- 22
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 3 ][ 6 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 2 ][ 6 ]; //  18 <- 19
assign fwd_data_in_o [ 2 ][ 7 ] = fwd_data_out_i [ 2 ][ 6 ]; //  19 -> 20
assign back_data_in_o[ 1 ][ 7 ] = back_data_out_i[ 1 ][ 6 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 1 ][ 6 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 6 ]; //  4 <- 5
assign fwd_data_in_o [ 0 ][ 7 ] = fwd_data_out_i [ 0 ][ 6 ]; //  5 -> 6
assign back_data_in_o[ 3 ][ 6 ] = back_data_out_i[ 3 ][ 5 ]; //  22 <- 23
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  23 -> 24
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  17 <- 18
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 2 ][ 5 ]; //  18 -> 19
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 1 ][ 5 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  23 <- 24
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  24 -> 25
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  16 <- 17
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  17 -> 18
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  10 -> 11
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  24 <- 25
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  25 -> 26
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  25 <- 26
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  26 -> 27
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  14 <- 15
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  11 <- 12
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  12 -> 13
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  26 <- 27
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 3 ][ 1 ]; //  27 -> 28
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  13 <- 14
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  13 -> 14
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  31 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 3 ][ 0 ]; //  27 <- 28
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  28 <- 29
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  29 -> 30
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  29 <- 30
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  30 -> 31
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  30 <- 31
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  31 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,  7,
  { b_lp ' (31) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4) , b_lp ' (5) , b_lp ' (6)     }, // x =  0
  { b_lp ' (30) , b_lp ' (13) , b_lp ' (12) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7)     }, // x =  1
  { b_lp ' (29) , b_lp ' (14) , b_lp ' (15) , b_lp ' (16) , b_lp ' (17) , b_lp ' (18) , b_lp ' (19) , b_lp ' (20)     }, // x =  2
  { b_lp ' (28) , b_lp ' (27) , b_lp ' (26) , b_lp ' (25) , b_lp ' (24) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21)     } // x =  3
 };
end
if (x_max_p == 6  && y_max_p == 2 )
begin
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 5 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 5 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  1 <- 2
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  2 -> 3
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  0 <- 1
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  11 <- 0
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 5 ][ 0 ]; //  5 <- 6
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  6 -> 7
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  6 <- 7
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  7 -> 8
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  8 -> 9
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  9 -> 10
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  9 <- 10
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  10 <- 11
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  11 -> 0
 assign id_o =
 {
// y =  0,  1,
  { b_lp ' (11) , b_lp ' (0)     }, // x =  0
  { b_lp ' (10) , b_lp ' (1)     }, // x =  1
  { b_lp ' (9) , b_lp ' (2)     }, // x =  2
  { b_lp ' (8) , b_lp ' (3)     }, // x =  3
  { b_lp ' (7) , b_lp ' (4)     }, // x =  4
  { b_lp ' (6) , b_lp ' (5)     } // x =  5
 };
end
if (x_max_p == 6  && y_max_p == 3 )
begin
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 5 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 4 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  5 <- 6
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  4 <- 5
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 1 ][ 2 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  2 -> 3
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 5 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  17 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 5 ][ 0 ]; //  11 <- 12
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  12 -> 13
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  12 <- 13
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  13 -> 14
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  13 <- 14
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  14 -> 15
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  14 <- 15
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  15 -> 16
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  15 <- 16
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  16 <- 17
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  17 -> 0
 assign id_o =
 {
// y =  0,  1,  2,
  { b_lp ' (17) , b_lp ' (0) , b_lp ' (1)     }, // x =  0
  { b_lp ' (16) , b_lp ' (3) , b_lp ' (2)     }, // x =  1
  { b_lp ' (15) , b_lp ' (4) , b_lp ' (5)     }, // x =  2
  { b_lp ' (14) , b_lp ' (7) , b_lp ' (6)     }, // x =  3
  { b_lp ' (13) , b_lp ' (8) , b_lp ' (9)     }, // x =  4
  { b_lp ' (12) , b_lp ' (11) , b_lp ' (10)     } // x =  5
 };
end
if (x_max_p == 6  && y_max_p == 4 )
begin
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 5 ][ 3 ]; //  14 <- 15
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  15 -> 16
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 4 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  8 <- 9
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  9 -> 10
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  7 <- 8
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  15 <- 16
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  16 -> 17
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  6 <- 7
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  7 -> 8
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  16 <- 17
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 5 ][ 1 ]; //  17 -> 18
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  11 <- 12
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  12 -> 13
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  23 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 5 ][ 0 ]; //  17 <- 18
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  18 -> 19
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  18 <- 19
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  19 -> 20
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  19 <- 20
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  20 -> 21
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  20 <- 21
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  21 <- 22
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  22 -> 23
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  22 <- 23
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  23 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,
  { b_lp ' (23) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2)     }, // x =  0
  { b_lp ' (22) , b_lp ' (5) , b_lp ' (4) , b_lp ' (3)     }, // x =  1
  { b_lp ' (21) , b_lp ' (6) , b_lp ' (7) , b_lp ' (8)     }, // x =  2
  { b_lp ' (20) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9)     }, // x =  3
  { b_lp ' (19) , b_lp ' (12) , b_lp ' (13) , b_lp ' (14)     }, // x =  4
  { b_lp ' (18) , b_lp ' (17) , b_lp ' (16) , b_lp ' (15)     } // x =  5
 };
end
if (x_max_p == 6  && y_max_p == 5 )
begin
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 5 ][ 4 ]; //  19 <- 20
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 5 ][ 4 ]; //  20 -> 21
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 4 ][ 4 ]; //  18 <- 19
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 4 ][ 4 ]; //  19 -> 20
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 3 ][ 4 ]; //  11 <- 12
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  12 -> 13
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  10 <- 11
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 2 ][ 4 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 1 ][ 4 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 5 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  17 <- 18
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 4 ][ 3 ]; //  18 -> 19
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  12 <- 13
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  13 -> 14
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  9 <- 10
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  21 <- 22
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  22 -> 23
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  16 <- 17
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  17 -> 18
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  13 <- 14
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  22 <- 23
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 5 ][ 1 ]; //  23 -> 24
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  15 <- 16
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  16 -> 17
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  14 <- 15
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  29 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 5 ][ 0 ]; //  23 <- 24
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  24 -> 25
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  24 <- 25
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  25 -> 26
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  25 <- 26
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  26 -> 27
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  26 <- 27
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  27 -> 28
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  27 <- 28
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  28 -> 29
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  28 <- 29
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  29 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,
  { b_lp ' (29) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3)     }, // x =  0
  { b_lp ' (28) , b_lp ' (7) , b_lp ' (6) , b_lp ' (5) , b_lp ' (4)     }, // x =  1
  { b_lp ' (27) , b_lp ' (8) , b_lp ' (9) , b_lp ' (10) , b_lp ' (11)     }, // x =  2
  { b_lp ' (26) , b_lp ' (15) , b_lp ' (14) , b_lp ' (13) , b_lp ' (12)     }, // x =  3
  { b_lp ' (25) , b_lp ' (16) , b_lp ' (17) , b_lp ' (18) , b_lp ' (19)     }, // x =  4
  { b_lp ' (24) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21) , b_lp ' (20)     } // x =  5
 };
end
if (x_max_p == 6  && y_max_p == 6 )
begin
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 5 ][ 5 ]; //  24 <- 25
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 5 ][ 5 ]; //  25 -> 26
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 4 ][ 5 ]; //  23 <- 24
assign fwd_data_in_o [ 5 ][ 5 ] = fwd_data_out_i [ 4 ][ 5 ]; //  24 -> 25
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 3 ][ 5 ]; //  14 <- 15
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  15 -> 16
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  13 <- 14
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  14 -> 15
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 5 ][ 5 ] = back_data_out_i[ 5 ][ 4 ]; //  25 <- 26
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 5 ][ 4 ]; //  26 -> 27
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 4 ][ 4 ]; //  22 <- 23
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 4 ][ 4 ]; //  23 -> 24
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  15 <- 16
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  16 -> 17
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 5 ][ 3 ]; //  26 <- 27
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  27 -> 28
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  21 <- 22
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 4 ][ 3 ]; //  22 -> 23
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  16 <- 17
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  17 -> 18
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  12 -> 13
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  27 <- 28
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  28 -> 29
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  20 <- 21
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  21 -> 22
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  17 <- 18
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  18 -> 19
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  10 <- 11
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  11 -> 12
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  28 <- 29
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 5 ][ 1 ]; //  29 -> 30
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  19 <- 20
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  20 -> 21
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  18 <- 19
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  19 -> 20
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  9 <- 10
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  35 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 5 ][ 0 ]; //  29 <- 30
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  30 -> 31
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  30 <- 31
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  31 -> 32
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  31 <- 32
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  32 -> 33
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  32 <- 33
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  33 -> 34
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  33 <- 34
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  34 -> 35
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  34 <- 35
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  35 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,
  { b_lp ' (35) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4)     }, // x =  0
  { b_lp ' (34) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7) , b_lp ' (6) , b_lp ' (5)     }, // x =  1
  { b_lp ' (33) , b_lp ' (10) , b_lp ' (11) , b_lp ' (12) , b_lp ' (13) , b_lp ' (14)     }, // x =  2
  { b_lp ' (32) , b_lp ' (19) , b_lp ' (18) , b_lp ' (17) , b_lp ' (16) , b_lp ' (15)     }, // x =  3
  { b_lp ' (31) , b_lp ' (20) , b_lp ' (21) , b_lp ' (22) , b_lp ' (23) , b_lp ' (24)     }, // x =  4
  { b_lp ' (30) , b_lp ' (29) , b_lp ' (28) , b_lp ' (27) , b_lp ' (26) , b_lp ' (25)     } // x =  5
 };
end
if (x_max_p == 6  && y_max_p == 7 )
begin
assign back_data_in_o[ 4 ][ 6 ] = back_data_out_i[ 5 ][ 6 ]; //  29 <- 30
assign fwd_data_in_o [ 5 ][ 5 ] = fwd_data_out_i [ 5 ][ 6 ]; //  30 -> 31
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 4 ][ 6 ]; //  28 <- 29
assign fwd_data_in_o [ 5 ][ 6 ] = fwd_data_out_i [ 4 ][ 6 ]; //  29 -> 30
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 3 ][ 6 ]; //  17 <- 18
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 3 ][ 6 ]; //  18 -> 19
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 2 ][ 6 ]; //  16 <- 17
assign fwd_data_in_o [ 3 ][ 6 ] = fwd_data_out_i [ 2 ][ 6 ]; //  17 -> 18
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 1 ][ 6 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 1 ][ 6 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 6 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 0 ][ 6 ]; //  5 -> 6
assign back_data_in_o[ 5 ][ 6 ] = back_data_out_i[ 5 ][ 5 ]; //  30 <- 31
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 5 ][ 5 ]; //  31 -> 32
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 4 ][ 5 ]; //  27 <- 28
assign fwd_data_in_o [ 4 ][ 6 ] = fwd_data_out_i [ 4 ][ 5 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 6 ] = back_data_out_i[ 3 ][ 5 ]; //  18 <- 19
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  19 -> 20
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 2 ][ 5 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 1 ][ 5 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 5 ][ 5 ] = back_data_out_i[ 5 ][ 4 ]; //  31 <- 32
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 5 ][ 4 ]; //  32 -> 33
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 4 ][ 4 ]; //  26 <- 27
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 4 ][ 4 ]; //  27 -> 28
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  20 -> 21
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  14 <- 15
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 5 ][ 3 ]; //  32 <- 33
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  33 -> 34
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  25 <- 26
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 4 ][ 3 ]; //  26 -> 27
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  33 <- 34
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  34 -> 35
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  24 <- 25
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  25 -> 26
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  21 <- 22
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  34 <- 35
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 5 ][ 1 ]; //  35 -> 36
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  23 <- 24
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  24 -> 25
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  22 <- 23
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  23 -> 24
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  12 -> 13
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  41 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 5 ][ 0 ]; //  35 <- 36
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  36 -> 37
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  36 <- 37
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  37 -> 38
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  37 <- 38
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  38 -> 39
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  38 <- 39
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  39 -> 40
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  39 <- 40
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  40 -> 41
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  40 <- 41
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  41 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,
  { b_lp ' (41) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4) , b_lp ' (5)     }, // x =  0
  { b_lp ' (40) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7) , b_lp ' (6)     }, // x =  1
  { b_lp ' (39) , b_lp ' (12) , b_lp ' (13) , b_lp ' (14) , b_lp ' (15) , b_lp ' (16) , b_lp ' (17)     }, // x =  2
  { b_lp ' (38) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21) , b_lp ' (20) , b_lp ' (19) , b_lp ' (18)     }, // x =  3
  { b_lp ' (37) , b_lp ' (24) , b_lp ' (25) , b_lp ' (26) , b_lp ' (27) , b_lp ' (28) , b_lp ' (29)     }, // x =  4
  { b_lp ' (36) , b_lp ' (35) , b_lp ' (34) , b_lp ' (33) , b_lp ' (32) , b_lp ' (31) , b_lp ' (30)     } // x =  5
 };
end
if (x_max_p == 6  && y_max_p == 8 )
begin
assign back_data_in_o[ 4 ][ 7 ] = back_data_out_i[ 5 ][ 7 ]; //  34 <- 35
assign fwd_data_in_o [ 5 ][ 6 ] = fwd_data_out_i [ 5 ][ 7 ]; //  35 -> 36
assign back_data_in_o[ 4 ][ 6 ] = back_data_out_i[ 4 ][ 7 ]; //  33 <- 34
assign fwd_data_in_o [ 5 ][ 7 ] = fwd_data_out_i [ 4 ][ 7 ]; //  34 -> 35
assign back_data_in_o[ 2 ][ 7 ] = back_data_out_i[ 3 ][ 7 ]; //  20 <- 21
assign fwd_data_in_o [ 3 ][ 6 ] = fwd_data_out_i [ 3 ][ 7 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 2 ][ 7 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 7 ] = fwd_data_out_i [ 2 ][ 7 ]; //  20 -> 21
assign back_data_in_o[ 0 ][ 7 ] = back_data_out_i[ 1 ][ 7 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 1 ][ 7 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 0 ][ 7 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 7 ] = fwd_data_out_i [ 0 ][ 7 ]; //  6 -> 7
assign back_data_in_o[ 5 ][ 7 ] = back_data_out_i[ 5 ][ 6 ]; //  35 <- 36
assign fwd_data_in_o [ 5 ][ 5 ] = fwd_data_out_i [ 5 ][ 6 ]; //  36 -> 37
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 4 ][ 6 ]; //  32 <- 33
assign fwd_data_in_o [ 4 ][ 7 ] = fwd_data_out_i [ 4 ][ 6 ]; //  33 -> 34
assign back_data_in_o[ 3 ][ 7 ] = back_data_out_i[ 3 ][ 6 ]; //  21 <- 22
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 3 ][ 6 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 2 ][ 6 ]; //  18 <- 19
assign fwd_data_in_o [ 2 ][ 7 ] = fwd_data_out_i [ 2 ][ 6 ]; //  19 -> 20
assign back_data_in_o[ 1 ][ 7 ] = back_data_out_i[ 1 ][ 6 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 1 ][ 6 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 6 ]; //  4 <- 5
assign fwd_data_in_o [ 0 ][ 7 ] = fwd_data_out_i [ 0 ][ 6 ]; //  5 -> 6
assign back_data_in_o[ 5 ][ 6 ] = back_data_out_i[ 5 ][ 5 ]; //  36 <- 37
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 5 ][ 5 ]; //  37 -> 38
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 4 ][ 5 ]; //  31 <- 32
assign fwd_data_in_o [ 4 ][ 6 ] = fwd_data_out_i [ 4 ][ 5 ]; //  32 -> 33
assign back_data_in_o[ 3 ][ 6 ] = back_data_out_i[ 3 ][ 5 ]; //  22 <- 23
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  23 -> 24
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  17 <- 18
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 2 ][ 5 ]; //  18 -> 19
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 1 ][ 5 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 5 ][ 5 ] = back_data_out_i[ 5 ][ 4 ]; //  37 <- 38
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 5 ][ 4 ]; //  38 -> 39
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 4 ][ 4 ]; //  30 <- 31
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 4 ][ 4 ]; //  31 -> 32
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  23 <- 24
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  24 -> 25
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  16 <- 17
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  17 -> 18
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  10 -> 11
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 5 ][ 3 ]; //  38 <- 39
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  39 -> 40
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  29 <- 30
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 4 ][ 3 ]; //  30 -> 31
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  24 <- 25
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  25 -> 26
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  39 <- 40
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  40 -> 41
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  28 <- 29
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  29 -> 30
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  25 <- 26
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  26 -> 27
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  14 <- 15
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  11 <- 12
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  12 -> 13
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  40 <- 41
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 5 ][ 1 ]; //  41 -> 42
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  27 <- 28
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  26 <- 27
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  27 -> 28
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  13 <- 14
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  13 -> 14
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  47 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 5 ][ 0 ]; //  41 <- 42
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  42 -> 43
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  42 <- 43
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  43 -> 44
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  43 <- 44
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  44 -> 45
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  44 <- 45
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  45 -> 46
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  45 <- 46
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  46 -> 47
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  46 <- 47
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  47 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,  7,
  { b_lp ' (47) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4) , b_lp ' (5) , b_lp ' (6)     }, // x =  0
  { b_lp ' (46) , b_lp ' (13) , b_lp ' (12) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7)     }, // x =  1
  { b_lp ' (45) , b_lp ' (14) , b_lp ' (15) , b_lp ' (16) , b_lp ' (17) , b_lp ' (18) , b_lp ' (19) , b_lp ' (20)     }, // x =  2
  { b_lp ' (44) , b_lp ' (27) , b_lp ' (26) , b_lp ' (25) , b_lp ' (24) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21)     }, // x =  3
  { b_lp ' (43) , b_lp ' (28) , b_lp ' (29) , b_lp ' (30) , b_lp ' (31) , b_lp ' (32) , b_lp ' (33) , b_lp ' (34)     }, // x =  4
  { b_lp ' (42) , b_lp ' (41) , b_lp ' (40) , b_lp ' (39) , b_lp ' (38) , b_lp ' (37) , b_lp ' (36) , b_lp ' (35)     } // x =  5
 };
end
if (x_max_p == 8  && y_max_p == 2 )
begin
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 7 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 7 ][ 0 ] = fwd_data_out_i [ 7 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 6 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 7 ][ 1 ] = fwd_data_out_i [ 6 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 5 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  1 <- 2
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  2 -> 3
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  0 <- 1
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  15 <- 0
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 7 ][ 1 ] = back_data_out_i[ 7 ][ 0 ]; //  7 <- 8
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 7 ][ 0 ]; //  8 -> 9
assign back_data_in_o[ 7 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  8 <- 9
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 6 ][ 0 ]; //  9 -> 10
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  9 <- 10
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  10 -> 11
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  10 <- 11
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  11 -> 12
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  12 -> 13
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  12 <- 13
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  13 -> 14
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  13 <- 14
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  14 <- 15
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  15 -> 0
 assign id_o =
 {
// y =  0,  1,
  { b_lp ' (15) , b_lp ' (0)     }, // x =  0
  { b_lp ' (14) , b_lp ' (1)     }, // x =  1
  { b_lp ' (13) , b_lp ' (2)     }, // x =  2
  { b_lp ' (12) , b_lp ' (3)     }, // x =  3
  { b_lp ' (11) , b_lp ' (4)     }, // x =  4
  { b_lp ' (10) , b_lp ' (5)     }, // x =  5
  { b_lp ' (9) , b_lp ' (6)     }, // x =  6
  { b_lp ' (8) , b_lp ' (7)     } // x =  7
 };
end
if (x_max_p == 8  && y_max_p == 3 )
begin
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 7 ][ 2 ]; //  13 <- 14
assign fwd_data_in_o [ 7 ][ 1 ] = fwd_data_out_i [ 7 ][ 2 ]; //  14 -> 15
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 6 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 7 ][ 2 ] = fwd_data_out_i [ 6 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 5 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 4 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  5 <- 6
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  4 <- 5
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 1 ][ 2 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  2 -> 3
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 7 ][ 2 ] = back_data_out_i[ 7 ][ 1 ]; //  14 <- 15
assign fwd_data_in_o [ 7 ][ 0 ] = fwd_data_out_i [ 7 ][ 1 ]; //  15 -> 16
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 6 ][ 1 ]; //  11 <- 12
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 6 ][ 1 ]; //  12 -> 13
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  23 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 7 ][ 1 ] = back_data_out_i[ 7 ][ 0 ]; //  15 <- 16
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 7 ][ 0 ]; //  16 -> 17
assign back_data_in_o[ 7 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  16 <- 17
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 6 ][ 0 ]; //  17 -> 18
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  17 <- 18
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  18 -> 19
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  18 <- 19
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  19 -> 20
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  19 <- 20
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  20 -> 21
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  20 <- 21
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  21 <- 22
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  22 -> 23
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  22 <- 23
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  23 -> 0
 assign id_o =
 {
// y =  0,  1,  2,
  { b_lp ' (23) , b_lp ' (0) , b_lp ' (1)     }, // x =  0
  { b_lp ' (22) , b_lp ' (3) , b_lp ' (2)     }, // x =  1
  { b_lp ' (21) , b_lp ' (4) , b_lp ' (5)     }, // x =  2
  { b_lp ' (20) , b_lp ' (7) , b_lp ' (6)     }, // x =  3
  { b_lp ' (19) , b_lp ' (8) , b_lp ' (9)     }, // x =  4
  { b_lp ' (18) , b_lp ' (11) , b_lp ' (10)     }, // x =  5
  { b_lp ' (17) , b_lp ' (12) , b_lp ' (13)     }, // x =  6
  { b_lp ' (16) , b_lp ' (15) , b_lp ' (14)     } // x =  7
 };
end
if (x_max_p == 8  && y_max_p == 4 )
begin
assign back_data_in_o[ 6 ][ 3 ] = back_data_out_i[ 7 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 7 ][ 2 ] = fwd_data_out_i [ 7 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 6 ][ 3 ]; //  19 <- 20
assign fwd_data_in_o [ 7 ][ 3 ] = fwd_data_out_i [ 6 ][ 3 ]; //  20 -> 21
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 5 ][ 3 ]; //  14 <- 15
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  15 -> 16
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 4 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  8 <- 9
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  9 -> 10
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  7 <- 8
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 7 ][ 3 ] = back_data_out_i[ 7 ][ 2 ]; //  21 <- 22
assign fwd_data_in_o [ 7 ][ 1 ] = fwd_data_out_i [ 7 ][ 2 ]; //  22 -> 23
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 6 ][ 2 ]; //  18 <- 19
assign fwd_data_in_o [ 6 ][ 3 ] = fwd_data_out_i [ 6 ][ 2 ]; //  19 -> 20
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  15 <- 16
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  16 -> 17
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  6 <- 7
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  7 -> 8
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 7 ][ 2 ] = back_data_out_i[ 7 ][ 1 ]; //  22 <- 23
assign fwd_data_in_o [ 7 ][ 0 ] = fwd_data_out_i [ 7 ][ 1 ]; //  23 -> 24
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 6 ][ 1 ]; //  17 <- 18
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 6 ][ 1 ]; //  18 -> 19
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  16 <- 17
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  17 -> 18
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  11 <- 12
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  12 -> 13
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  31 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 7 ][ 1 ] = back_data_out_i[ 7 ][ 0 ]; //  23 <- 24
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 7 ][ 0 ]; //  24 -> 25
assign back_data_in_o[ 7 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  24 <- 25
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 6 ][ 0 ]; //  25 -> 26
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  25 <- 26
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  26 -> 27
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  26 <- 27
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  27 -> 28
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  27 <- 28
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  28 <- 29
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  29 -> 30
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  29 <- 30
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  30 -> 31
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  30 <- 31
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  31 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,
  { b_lp ' (31) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2)     }, // x =  0
  { b_lp ' (30) , b_lp ' (5) , b_lp ' (4) , b_lp ' (3)     }, // x =  1
  { b_lp ' (29) , b_lp ' (6) , b_lp ' (7) , b_lp ' (8)     }, // x =  2
  { b_lp ' (28) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9)     }, // x =  3
  { b_lp ' (27) , b_lp ' (12) , b_lp ' (13) , b_lp ' (14)     }, // x =  4
  { b_lp ' (26) , b_lp ' (17) , b_lp ' (16) , b_lp ' (15)     }, // x =  5
  { b_lp ' (25) , b_lp ' (18) , b_lp ' (19) , b_lp ' (20)     }, // x =  6
  { b_lp ' (24) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21)     } // x =  7
 };
end
if (x_max_p == 8  && y_max_p == 5 )
begin
assign back_data_in_o[ 6 ][ 4 ] = back_data_out_i[ 7 ][ 4 ]; //  27 <- 28
assign fwd_data_in_o [ 7 ][ 3 ] = fwd_data_out_i [ 7 ][ 4 ]; //  28 -> 29
assign back_data_in_o[ 6 ][ 3 ] = back_data_out_i[ 6 ][ 4 ]; //  26 <- 27
assign fwd_data_in_o [ 7 ][ 4 ] = fwd_data_out_i [ 6 ][ 4 ]; //  27 -> 28
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 5 ][ 4 ]; //  19 <- 20
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 5 ][ 4 ]; //  20 -> 21
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 4 ][ 4 ]; //  18 <- 19
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 4 ][ 4 ]; //  19 -> 20
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 3 ][ 4 ]; //  11 <- 12
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  12 -> 13
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  10 <- 11
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 2 ][ 4 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 1 ][ 4 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 7 ][ 4 ] = back_data_out_i[ 7 ][ 3 ]; //  28 <- 29
assign fwd_data_in_o [ 7 ][ 2 ] = fwd_data_out_i [ 7 ][ 3 ]; //  29 -> 30
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 6 ][ 3 ]; //  25 <- 26
assign fwd_data_in_o [ 6 ][ 4 ] = fwd_data_out_i [ 6 ][ 3 ]; //  26 -> 27
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 5 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  17 <- 18
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 4 ][ 3 ]; //  18 -> 19
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  12 <- 13
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  13 -> 14
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  9 <- 10
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 7 ][ 3 ] = back_data_out_i[ 7 ][ 2 ]; //  29 <- 30
assign fwd_data_in_o [ 7 ][ 1 ] = fwd_data_out_i [ 7 ][ 2 ]; //  30 -> 31
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 6 ][ 2 ]; //  24 <- 25
assign fwd_data_in_o [ 6 ][ 3 ] = fwd_data_out_i [ 6 ][ 2 ]; //  25 -> 26
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  21 <- 22
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  22 -> 23
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  16 <- 17
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  17 -> 18
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  13 <- 14
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 7 ][ 2 ] = back_data_out_i[ 7 ][ 1 ]; //  30 <- 31
assign fwd_data_in_o [ 7 ][ 0 ] = fwd_data_out_i [ 7 ][ 1 ]; //  31 -> 32
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 6 ][ 1 ]; //  23 <- 24
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 6 ][ 1 ]; //  24 -> 25
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  22 <- 23
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  23 -> 24
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  15 <- 16
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  16 -> 17
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  14 <- 15
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  39 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 7 ][ 1 ] = back_data_out_i[ 7 ][ 0 ]; //  31 <- 32
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 7 ][ 0 ]; //  32 -> 33
assign back_data_in_o[ 7 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  32 <- 33
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 6 ][ 0 ]; //  33 -> 34
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  33 <- 34
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  34 -> 35
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  34 <- 35
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  35 -> 36
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  35 <- 36
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  36 -> 37
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  36 <- 37
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  37 -> 38
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  37 <- 38
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  38 -> 39
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  38 <- 39
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  39 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,
  { b_lp ' (39) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3)     }, // x =  0
  { b_lp ' (38) , b_lp ' (7) , b_lp ' (6) , b_lp ' (5) , b_lp ' (4)     }, // x =  1
  { b_lp ' (37) , b_lp ' (8) , b_lp ' (9) , b_lp ' (10) , b_lp ' (11)     }, // x =  2
  { b_lp ' (36) , b_lp ' (15) , b_lp ' (14) , b_lp ' (13) , b_lp ' (12)     }, // x =  3
  { b_lp ' (35) , b_lp ' (16) , b_lp ' (17) , b_lp ' (18) , b_lp ' (19)     }, // x =  4
  { b_lp ' (34) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21) , b_lp ' (20)     }, // x =  5
  { b_lp ' (33) , b_lp ' (24) , b_lp ' (25) , b_lp ' (26) , b_lp ' (27)     }, // x =  6
  { b_lp ' (32) , b_lp ' (31) , b_lp ' (30) , b_lp ' (29) , b_lp ' (28)     } // x =  7
 };
end
if (x_max_p == 8  && y_max_p == 6 )
begin
assign back_data_in_o[ 6 ][ 5 ] = back_data_out_i[ 7 ][ 5 ]; //  34 <- 35
assign fwd_data_in_o [ 7 ][ 4 ] = fwd_data_out_i [ 7 ][ 5 ]; //  35 -> 36
assign back_data_in_o[ 6 ][ 4 ] = back_data_out_i[ 6 ][ 5 ]; //  33 <- 34
assign fwd_data_in_o [ 7 ][ 5 ] = fwd_data_out_i [ 6 ][ 5 ]; //  34 -> 35
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 5 ][ 5 ]; //  24 <- 25
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 5 ][ 5 ]; //  25 -> 26
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 4 ][ 5 ]; //  23 <- 24
assign fwd_data_in_o [ 5 ][ 5 ] = fwd_data_out_i [ 4 ][ 5 ]; //  24 -> 25
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 3 ][ 5 ]; //  14 <- 15
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  15 -> 16
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  13 <- 14
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  14 -> 15
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  5 -> 6
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 7 ][ 5 ] = back_data_out_i[ 7 ][ 4 ]; //  35 <- 36
assign fwd_data_in_o [ 7 ][ 3 ] = fwd_data_out_i [ 7 ][ 4 ]; //  36 -> 37
assign back_data_in_o[ 6 ][ 3 ] = back_data_out_i[ 6 ][ 4 ]; //  32 <- 33
assign fwd_data_in_o [ 6 ][ 5 ] = fwd_data_out_i [ 6 ][ 4 ]; //  33 -> 34
assign back_data_in_o[ 5 ][ 5 ] = back_data_out_i[ 5 ][ 4 ]; //  25 <- 26
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 5 ][ 4 ]; //  26 -> 27
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 4 ][ 4 ]; //  22 <- 23
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 4 ][ 4 ]; //  23 -> 24
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  15 <- 16
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  16 -> 17
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 7 ][ 4 ] = back_data_out_i[ 7 ][ 3 ]; //  36 <- 37
assign fwd_data_in_o [ 7 ][ 2 ] = fwd_data_out_i [ 7 ][ 3 ]; //  37 -> 38
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 6 ][ 3 ]; //  31 <- 32
assign fwd_data_in_o [ 6 ][ 4 ] = fwd_data_out_i [ 6 ][ 3 ]; //  32 -> 33
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 5 ][ 3 ]; //  26 <- 27
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  27 -> 28
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  21 <- 22
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 4 ][ 3 ]; //  22 -> 23
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  16 <- 17
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  17 -> 18
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  12 -> 13
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 7 ][ 3 ] = back_data_out_i[ 7 ][ 2 ]; //  37 <- 38
assign fwd_data_in_o [ 7 ][ 1 ] = fwd_data_out_i [ 7 ][ 2 ]; //  38 -> 39
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 6 ][ 2 ]; //  30 <- 31
assign fwd_data_in_o [ 6 ][ 3 ] = fwd_data_out_i [ 6 ][ 2 ]; //  31 -> 32
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  27 <- 28
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  28 -> 29
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  20 <- 21
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  21 -> 22
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  17 <- 18
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  18 -> 19
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  10 <- 11
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  11 -> 12
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 7 ][ 2 ] = back_data_out_i[ 7 ][ 1 ]; //  38 <- 39
assign fwd_data_in_o [ 7 ][ 0 ] = fwd_data_out_i [ 7 ][ 1 ]; //  39 -> 40
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 6 ][ 1 ]; //  29 <- 30
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 6 ][ 1 ]; //  30 -> 31
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  28 <- 29
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  29 -> 30
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  19 <- 20
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  20 -> 21
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  18 <- 19
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  19 -> 20
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  9 <- 10
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  47 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 7 ][ 1 ] = back_data_out_i[ 7 ][ 0 ]; //  39 <- 40
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 7 ][ 0 ]; //  40 -> 41
assign back_data_in_o[ 7 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  40 <- 41
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 6 ][ 0 ]; //  41 -> 42
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  41 <- 42
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  42 -> 43
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  42 <- 43
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  43 -> 44
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  43 <- 44
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  44 -> 45
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  44 <- 45
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  45 -> 46
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  45 <- 46
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  46 -> 47
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  46 <- 47
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  47 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,
  { b_lp ' (47) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4)     }, // x =  0
  { b_lp ' (46) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7) , b_lp ' (6) , b_lp ' (5)     }, // x =  1
  { b_lp ' (45) , b_lp ' (10) , b_lp ' (11) , b_lp ' (12) , b_lp ' (13) , b_lp ' (14)     }, // x =  2
  { b_lp ' (44) , b_lp ' (19) , b_lp ' (18) , b_lp ' (17) , b_lp ' (16) , b_lp ' (15)     }, // x =  3
  { b_lp ' (43) , b_lp ' (20) , b_lp ' (21) , b_lp ' (22) , b_lp ' (23) , b_lp ' (24)     }, // x =  4
  { b_lp ' (42) , b_lp ' (29) , b_lp ' (28) , b_lp ' (27) , b_lp ' (26) , b_lp ' (25)     }, // x =  5
  { b_lp ' (41) , b_lp ' (30) , b_lp ' (31) , b_lp ' (32) , b_lp ' (33) , b_lp ' (34)     }, // x =  6
  { b_lp ' (40) , b_lp ' (39) , b_lp ' (38) , b_lp ' (37) , b_lp ' (36) , b_lp ' (35)     } // x =  7
 };
end
if (x_max_p == 8  && y_max_p == 7 )
begin
assign back_data_in_o[ 6 ][ 6 ] = back_data_out_i[ 7 ][ 6 ]; //  41 <- 42
assign fwd_data_in_o [ 7 ][ 5 ] = fwd_data_out_i [ 7 ][ 6 ]; //  42 -> 43
assign back_data_in_o[ 6 ][ 5 ] = back_data_out_i[ 6 ][ 6 ]; //  40 <- 41
assign fwd_data_in_o [ 7 ][ 6 ] = fwd_data_out_i [ 6 ][ 6 ]; //  41 -> 42
assign back_data_in_o[ 4 ][ 6 ] = back_data_out_i[ 5 ][ 6 ]; //  29 <- 30
assign fwd_data_in_o [ 5 ][ 5 ] = fwd_data_out_i [ 5 ][ 6 ]; //  30 -> 31
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 4 ][ 6 ]; //  28 <- 29
assign fwd_data_in_o [ 5 ][ 6 ] = fwd_data_out_i [ 4 ][ 6 ]; //  29 -> 30
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 3 ][ 6 ]; //  17 <- 18
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 3 ][ 6 ]; //  18 -> 19
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 2 ][ 6 ]; //  16 <- 17
assign fwd_data_in_o [ 3 ][ 6 ] = fwd_data_out_i [ 2 ][ 6 ]; //  17 -> 18
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 1 ][ 6 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 1 ][ 6 ]; //  6 -> 7
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 6 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 0 ][ 6 ]; //  5 -> 6
assign back_data_in_o[ 7 ][ 6 ] = back_data_out_i[ 7 ][ 5 ]; //  42 <- 43
assign fwd_data_in_o [ 7 ][ 4 ] = fwd_data_out_i [ 7 ][ 5 ]; //  43 -> 44
assign back_data_in_o[ 6 ][ 4 ] = back_data_out_i[ 6 ][ 5 ]; //  39 <- 40
assign fwd_data_in_o [ 6 ][ 6 ] = fwd_data_out_i [ 6 ][ 5 ]; //  40 -> 41
assign back_data_in_o[ 5 ][ 6 ] = back_data_out_i[ 5 ][ 5 ]; //  30 <- 31
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 5 ][ 5 ]; //  31 -> 32
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 4 ][ 5 ]; //  27 <- 28
assign fwd_data_in_o [ 4 ][ 6 ] = fwd_data_out_i [ 4 ][ 5 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 6 ] = back_data_out_i[ 3 ][ 5 ]; //  18 <- 19
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  19 -> 20
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 2 ][ 5 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 1 ][ 5 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 7 ][ 5 ] = back_data_out_i[ 7 ][ 4 ]; //  43 <- 44
assign fwd_data_in_o [ 7 ][ 3 ] = fwd_data_out_i [ 7 ][ 4 ]; //  44 -> 45
assign back_data_in_o[ 6 ][ 3 ] = back_data_out_i[ 6 ][ 4 ]; //  38 <- 39
assign fwd_data_in_o [ 6 ][ 5 ] = fwd_data_out_i [ 6 ][ 4 ]; //  39 -> 40
assign back_data_in_o[ 5 ][ 5 ] = back_data_out_i[ 5 ][ 4 ]; //  31 <- 32
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 5 ][ 4 ]; //  32 -> 33
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 4 ][ 4 ]; //  26 <- 27
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 4 ][ 4 ]; //  27 -> 28
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  20 -> 21
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  14 <- 15
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 7 ][ 4 ] = back_data_out_i[ 7 ][ 3 ]; //  44 <- 45
assign fwd_data_in_o [ 7 ][ 2 ] = fwd_data_out_i [ 7 ][ 3 ]; //  45 -> 46
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 6 ][ 3 ]; //  37 <- 38
assign fwd_data_in_o [ 6 ][ 4 ] = fwd_data_out_i [ 6 ][ 3 ]; //  38 -> 39
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 5 ][ 3 ]; //  32 <- 33
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  33 -> 34
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  25 <- 26
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 4 ][ 3 ]; //  26 -> 27
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 7 ][ 3 ] = back_data_out_i[ 7 ][ 2 ]; //  45 <- 46
assign fwd_data_in_o [ 7 ][ 1 ] = fwd_data_out_i [ 7 ][ 2 ]; //  46 -> 47
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 6 ][ 2 ]; //  36 <- 37
assign fwd_data_in_o [ 6 ][ 3 ] = fwd_data_out_i [ 6 ][ 2 ]; //  37 -> 38
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  33 <- 34
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  34 -> 35
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  24 <- 25
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  25 -> 26
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  21 <- 22
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 7 ][ 2 ] = back_data_out_i[ 7 ][ 1 ]; //  46 <- 47
assign fwd_data_in_o [ 7 ][ 0 ] = fwd_data_out_i [ 7 ][ 1 ]; //  47 -> 48
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 6 ][ 1 ]; //  35 <- 36
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 6 ][ 1 ]; //  36 -> 37
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  34 <- 35
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  35 -> 36
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  23 <- 24
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  24 -> 25
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  22 <- 23
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  23 -> 24
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  12 -> 13
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  55 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 7 ][ 1 ] = back_data_out_i[ 7 ][ 0 ]; //  47 <- 48
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 7 ][ 0 ]; //  48 -> 49
assign back_data_in_o[ 7 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  48 <- 49
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 6 ][ 0 ]; //  49 -> 50
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  49 <- 50
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  50 -> 51
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  50 <- 51
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  51 -> 52
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  51 <- 52
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  52 -> 53
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  52 <- 53
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  53 -> 54
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  53 <- 54
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  54 -> 55
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  54 <- 55
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  55 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,
  { b_lp ' (55) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4) , b_lp ' (5)     }, // x =  0
  { b_lp ' (54) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7) , b_lp ' (6)     }, // x =  1
  { b_lp ' (53) , b_lp ' (12) , b_lp ' (13) , b_lp ' (14) , b_lp ' (15) , b_lp ' (16) , b_lp ' (17)     }, // x =  2
  { b_lp ' (52) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21) , b_lp ' (20) , b_lp ' (19) , b_lp ' (18)     }, // x =  3
  { b_lp ' (51) , b_lp ' (24) , b_lp ' (25) , b_lp ' (26) , b_lp ' (27) , b_lp ' (28) , b_lp ' (29)     }, // x =  4
  { b_lp ' (50) , b_lp ' (35) , b_lp ' (34) , b_lp ' (33) , b_lp ' (32) , b_lp ' (31) , b_lp ' (30)     }, // x =  5
  { b_lp ' (49) , b_lp ' (36) , b_lp ' (37) , b_lp ' (38) , b_lp ' (39) , b_lp ' (40) , b_lp ' (41)     }, // x =  6
  { b_lp ' (48) , b_lp ' (47) , b_lp ' (46) , b_lp ' (45) , b_lp ' (44) , b_lp ' (43) , b_lp ' (42)     } // x =  7
 };
end
if (x_max_p == 8  && y_max_p == 8 )
begin
assign back_data_in_o[ 6 ][ 7 ] = back_data_out_i[ 7 ][ 7 ]; //  48 <- 49
assign fwd_data_in_o [ 7 ][ 6 ] = fwd_data_out_i [ 7 ][ 7 ]; //  49 -> 50
assign back_data_in_o[ 6 ][ 6 ] = back_data_out_i[ 6 ][ 7 ]; //  47 <- 48
assign fwd_data_in_o [ 7 ][ 7 ] = fwd_data_out_i [ 6 ][ 7 ]; //  48 -> 49
assign back_data_in_o[ 4 ][ 7 ] = back_data_out_i[ 5 ][ 7 ]; //  34 <- 35
assign fwd_data_in_o [ 5 ][ 6 ] = fwd_data_out_i [ 5 ][ 7 ]; //  35 -> 36
assign back_data_in_o[ 4 ][ 6 ] = back_data_out_i[ 4 ][ 7 ]; //  33 <- 34
assign fwd_data_in_o [ 5 ][ 7 ] = fwd_data_out_i [ 4 ][ 7 ]; //  34 -> 35
assign back_data_in_o[ 2 ][ 7 ] = back_data_out_i[ 3 ][ 7 ]; //  20 <- 21
assign fwd_data_in_o [ 3 ][ 6 ] = fwd_data_out_i [ 3 ][ 7 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 2 ][ 7 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 7 ] = fwd_data_out_i [ 2 ][ 7 ]; //  20 -> 21
assign back_data_in_o[ 0 ][ 7 ] = back_data_out_i[ 1 ][ 7 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 1 ][ 7 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 0 ][ 7 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 7 ] = fwd_data_out_i [ 0 ][ 7 ]; //  6 -> 7
assign back_data_in_o[ 7 ][ 7 ] = back_data_out_i[ 7 ][ 6 ]; //  49 <- 50
assign fwd_data_in_o [ 7 ][ 5 ] = fwd_data_out_i [ 7 ][ 6 ]; //  50 -> 51
assign back_data_in_o[ 6 ][ 5 ] = back_data_out_i[ 6 ][ 6 ]; //  46 <- 47
assign fwd_data_in_o [ 6 ][ 7 ] = fwd_data_out_i [ 6 ][ 6 ]; //  47 -> 48
assign back_data_in_o[ 5 ][ 7 ] = back_data_out_i[ 5 ][ 6 ]; //  35 <- 36
assign fwd_data_in_o [ 5 ][ 5 ] = fwd_data_out_i [ 5 ][ 6 ]; //  36 -> 37
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 4 ][ 6 ]; //  32 <- 33
assign fwd_data_in_o [ 4 ][ 7 ] = fwd_data_out_i [ 4 ][ 6 ]; //  33 -> 34
assign back_data_in_o[ 3 ][ 7 ] = back_data_out_i[ 3 ][ 6 ]; //  21 <- 22
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 3 ][ 6 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 2 ][ 6 ]; //  18 <- 19
assign fwd_data_in_o [ 2 ][ 7 ] = fwd_data_out_i [ 2 ][ 6 ]; //  19 -> 20
assign back_data_in_o[ 1 ][ 7 ] = back_data_out_i[ 1 ][ 6 ]; //  7 <- 8
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 1 ][ 6 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 6 ]; //  4 <- 5
assign fwd_data_in_o [ 0 ][ 7 ] = fwd_data_out_i [ 0 ][ 6 ]; //  5 -> 6
assign back_data_in_o[ 7 ][ 6 ] = back_data_out_i[ 7 ][ 5 ]; //  50 <- 51
assign fwd_data_in_o [ 7 ][ 4 ] = fwd_data_out_i [ 7 ][ 5 ]; //  51 -> 52
assign back_data_in_o[ 6 ][ 4 ] = back_data_out_i[ 6 ][ 5 ]; //  45 <- 46
assign fwd_data_in_o [ 6 ][ 6 ] = fwd_data_out_i [ 6 ][ 5 ]; //  46 -> 47
assign back_data_in_o[ 5 ][ 6 ] = back_data_out_i[ 5 ][ 5 ]; //  36 <- 37
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 5 ][ 5 ]; //  37 -> 38
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 4 ][ 5 ]; //  31 <- 32
assign fwd_data_in_o [ 4 ][ 6 ] = fwd_data_out_i [ 4 ][ 5 ]; //  32 -> 33
assign back_data_in_o[ 3 ][ 6 ] = back_data_out_i[ 3 ][ 5 ]; //  22 <- 23
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 3 ][ 5 ]; //  23 -> 24
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  17 <- 18
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 2 ][ 5 ]; //  18 -> 19
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 1 ][ 5 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 5 ]; //  9 -> 10
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 5 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 5 ]; //  4 -> 5
assign back_data_in_o[ 7 ][ 5 ] = back_data_out_i[ 7 ][ 4 ]; //  51 <- 52
assign fwd_data_in_o [ 7 ][ 3 ] = fwd_data_out_i [ 7 ][ 4 ]; //  52 -> 53
assign back_data_in_o[ 6 ][ 3 ] = back_data_out_i[ 6 ][ 4 ]; //  44 <- 45
assign fwd_data_in_o [ 6 ][ 5 ] = fwd_data_out_i [ 6 ][ 4 ]; //  45 -> 46
assign back_data_in_o[ 5 ][ 5 ] = back_data_out_i[ 5 ][ 4 ]; //  37 <- 38
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 5 ][ 4 ]; //  38 -> 39
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 4 ][ 4 ]; //  30 <- 31
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 4 ][ 4 ]; //  31 -> 32
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 3 ][ 4 ]; //  23 <- 24
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 3 ][ 4 ]; //  24 -> 25
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 2 ][ 4 ]; //  16 <- 17
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  17 -> 18
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 4 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 1 ][ 4 ]; //  10 -> 11
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 4 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 4 ]; //  3 -> 4
assign back_data_in_o[ 7 ][ 4 ] = back_data_out_i[ 7 ][ 3 ]; //  52 <- 53
assign fwd_data_in_o [ 7 ][ 2 ] = fwd_data_out_i [ 7 ][ 3 ]; //  53 -> 54
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 6 ][ 3 ]; //  43 <- 44
assign fwd_data_in_o [ 6 ][ 4 ] = fwd_data_out_i [ 6 ][ 3 ]; //  44 -> 45
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 5 ][ 3 ]; //  38 <- 39
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 5 ][ 3 ]; //  39 -> 40
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  29 <- 30
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 4 ][ 3 ]; //  30 -> 31
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 3 ][ 3 ]; //  24 <- 25
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 3 ][ 3 ]; //  25 -> 26
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 2 ][ 3 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 1 ][ 3 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 3 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 3 ]; //  1 <- 2
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 3 ]; //  2 -> 3
assign back_data_in_o[ 7 ][ 3 ] = back_data_out_i[ 7 ][ 2 ]; //  53 <- 54
assign fwd_data_in_o [ 7 ][ 1 ] = fwd_data_out_i [ 7 ][ 2 ]; //  54 -> 55
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 6 ][ 2 ]; //  42 <- 43
assign fwd_data_in_o [ 6 ][ 3 ] = fwd_data_out_i [ 6 ][ 2 ]; //  43 -> 44
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 5 ][ 2 ]; //  39 <- 40
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 5 ][ 2 ]; //  40 -> 41
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 4 ][ 2 ]; //  28 <- 29
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  29 -> 30
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 3 ][ 2 ]; //  25 <- 26
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 3 ][ 2 ]; //  26 -> 27
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 2 ][ 2 ]; //  14 <- 15
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 2 ]; //  11 <- 12
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 1 ][ 2 ]; //  12 -> 13
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 2 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 2 ]; //  1 -> 2
assign back_data_in_o[ 7 ][ 2 ] = back_data_out_i[ 7 ][ 1 ]; //  54 <- 55
assign fwd_data_in_o [ 7 ][ 0 ] = fwd_data_out_i [ 7 ][ 1 ]; //  55 -> 56
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 6 ][ 1 ]; //  41 <- 42
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 6 ][ 1 ]; //  42 -> 43
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 5 ][ 1 ]; //  40 <- 41
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  41 -> 42
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  27 <- 28
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 4 ][ 1 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 3 ][ 1 ]; //  26 <- 27
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  27 -> 28
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  13 <- 14
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 2 ][ 1 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 1 ][ 1 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  13 -> 14
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  63 <- 0
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 1 ]; //  0 -> 1
assign back_data_in_o[ 7 ][ 1 ] = back_data_out_i[ 7 ][ 0 ]; //  55 <- 56
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 7 ][ 0 ]; //  56 -> 57
assign back_data_in_o[ 7 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  56 <- 57
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 6 ][ 0 ]; //  57 -> 58
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  57 <- 58
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  58 -> 59
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  58 <- 59
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  59 -> 60
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  59 <- 60
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  60 -> 61
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  60 <- 61
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  61 -> 62
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  61 <- 62
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  62 -> 63
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  62 <- 63
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  63 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,  7,
  { b_lp ' (63) , b_lp ' (0) , b_lp ' (1) , b_lp ' (2) , b_lp ' (3) , b_lp ' (4) , b_lp ' (5) , b_lp ' (6)     }, // x =  0
  { b_lp ' (62) , b_lp ' (13) , b_lp ' (12) , b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8) , b_lp ' (7)     }, // x =  1
  { b_lp ' (61) , b_lp ' (14) , b_lp ' (15) , b_lp ' (16) , b_lp ' (17) , b_lp ' (18) , b_lp ' (19) , b_lp ' (20)     }, // x =  2
  { b_lp ' (60) , b_lp ' (27) , b_lp ' (26) , b_lp ' (25) , b_lp ' (24) , b_lp ' (23) , b_lp ' (22) , b_lp ' (21)     }, // x =  3
  { b_lp ' (59) , b_lp ' (28) , b_lp ' (29) , b_lp ' (30) , b_lp ' (31) , b_lp ' (32) , b_lp ' (33) , b_lp ' (34)     }, // x =  4
  { b_lp ' (58) , b_lp ' (41) , b_lp ' (40) , b_lp ' (39) , b_lp ' (38) , b_lp ' (37) , b_lp ' (36) , b_lp ' (35)     }, // x =  5
  { b_lp ' (57) , b_lp ' (42) , b_lp ' (43) , b_lp ' (44) , b_lp ' (45) , b_lp ' (46) , b_lp ' (47) , b_lp ' (48)     }, // x =  6
  { b_lp ' (56) , b_lp ' (55) , b_lp ' (54) , b_lp ' (53) , b_lp ' (52) , b_lp ' (51) , b_lp ' (50) , b_lp ' (49)     } // x =  7
 };
end
if (x_max_p == 3  && y_max_p == 2 )
begin
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 2 ][ 1 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  2 -> 3
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 0 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  5 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  4 <- 5
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  5 -> 0
 assign id_o =
 {
// y =  0,  1,
  { b_lp ' (5) , b_lp ' (4)     }, // x =  0
  { b_lp ' (0) , b_lp ' (3)     }, // x =  1
  { b_lp ' (1) , b_lp ' (2)     } // x =  2
 };
end
if (x_max_p == 3  && y_max_p == 4 )
begin
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  6 <- 7
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 1 ][ 3 ]; //  7 -> 8
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 0 ][ 3 ]; //  7 <- 8
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  8 -> 9
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  5 -> 6
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  3 <- 4
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 2 ][ 1 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  2 -> 3
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  9 <- 10
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  11 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  11 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,
  { b_lp ' (11) , b_lp ' (10) , b_lp ' (9) , b_lp ' (8)     }, // x =  0
  { b_lp ' (0) , b_lp ' (3) , b_lp ' (4) , b_lp ' (7)     }, // x =  1
  { b_lp ' (1) , b_lp ' (2) , b_lp ' (5) , b_lp ' (6)     } // x =  2
 };
end
if (x_max_p == 3  && y_max_p == 6 )
begin
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  10 <- 11
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 1 ][ 5 ]; //  11 -> 12
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 0 ][ 5 ]; //  11 <- 12
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 5 ]; //  12 -> 13
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 2 ][ 4 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  9 -> 10
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 4 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 1 ][ 4 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 4 ]; //  12 <- 13
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 4 ]; //  13 -> 14
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 3 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  5 -> 6
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  3 <- 4
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  14 <- 15
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  15 -> 16
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 2 ][ 1 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  2 -> 3
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  15 <- 16
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  17 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  16 <- 17
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  17 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,
  { b_lp ' (17) , b_lp ' (16) , b_lp ' (15) , b_lp ' (14) , b_lp ' (13) , b_lp ' (12)     }, // x =  0
  { b_lp ' (0) , b_lp ' (3) , b_lp ' (4) , b_lp ' (7) , b_lp ' (8) , b_lp ' (11)     }, // x =  1
  { b_lp ' (1) , b_lp ' (2) , b_lp ' (5) , b_lp ' (6) , b_lp ' (9) , b_lp ' (10)     } // x =  2
 };
end
if (x_max_p == 3  && y_max_p == 8 )
begin
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 2 ][ 7 ]; //  13 <- 14
assign fwd_data_in_o [ 1 ][ 7 ] = fwd_data_out_i [ 2 ][ 7 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 7 ] = back_data_out_i[ 1 ][ 7 ]; //  14 <- 15
assign fwd_data_in_o [ 0 ][ 7 ] = fwd_data_out_i [ 1 ][ 7 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 7 ] = back_data_out_i[ 0 ][ 7 ]; //  15 <- 16
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 7 ]; //  16 -> 17
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 2 ][ 6 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 7 ] = fwd_data_out_i [ 2 ][ 6 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 6 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 1 ][ 6 ]; //  12 -> 13
assign back_data_in_o[ 0 ][ 7 ] = back_data_out_i[ 0 ][ 6 ]; //  16 <- 17
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 6 ]; //  17 -> 18
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 2 ][ 5 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 1 ][ 5 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 0 ][ 5 ]; //  17 <- 18
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 5 ]; //  18 -> 19
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 2 ][ 4 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 2 ][ 4 ]; //  9 -> 10
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 4 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 1 ][ 4 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 4 ]; //  18 <- 19
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 4 ]; //  19 -> 20
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 2 ][ 3 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 3 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 3 ]; //  19 <- 20
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  20 -> 21
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 2 ][ 2 ]; //  5 -> 6
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  3 <- 4
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  4 -> 5
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  20 <- 21
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  21 -> 22
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 2 ][ 1 ]; //  1 <- 2
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  2 -> 3
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  2 <- 3
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  3 -> 4
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  21 <- 22
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  22 -> 23
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  23 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  22 <- 23
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  23 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,  7,
  { b_lp ' (23) , b_lp ' (22) , b_lp ' (21) , b_lp ' (20) , b_lp ' (19) , b_lp ' (18) , b_lp ' (17) , b_lp ' (16)     }, // x =  0
  { b_lp ' (0) , b_lp ' (3) , b_lp ' (4) , b_lp ' (7) , b_lp ' (8) , b_lp ' (11) , b_lp ' (12) , b_lp ' (15)     }, // x =  1
  { b_lp ' (1) , b_lp ' (2) , b_lp ' (5) , b_lp ' (6) , b_lp ' (9) , b_lp ' (10) , b_lp ' (13) , b_lp ' (14)     } // x =  2
 };
end
if (x_max_p == 5  && y_max_p == 2 )
begin
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 4 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 0 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 4 ][ 0 ]; //  3 -> 4
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  9 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  8 <- 9
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  9 -> 0
 assign id_o =
 {
// y =  0,  1,
  { b_lp ' (9) , b_lp ' (8)     }, // x =  0
  { b_lp ' (0) , b_lp ' (7)     }, // x =  1
  { b_lp ' (1) , b_lp ' (6)     }, // x =  2
  { b_lp ' (2) , b_lp ' (5)     }, // x =  3
  { b_lp ' (3) , b_lp ' (4)     } // x =  4
 };
end
if (x_max_p == 5  && y_max_p == 4 )
begin
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  11 <- 12
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 4 ][ 3 ]; //  12 -> 13
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 3 ][ 3 ]; //  13 -> 14
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 2 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  14 <- 15
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 1 ][ 3 ]; //  15 -> 16
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 0 ][ 3 ]; //  15 <- 16
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  16 -> 17
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 4 ][ 2 ]; //  10 <- 11
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  11 -> 12
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 3 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  16 <- 17
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  17 -> 18
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 4 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  17 <- 18
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  18 -> 19
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 4 ][ 0 ]; //  3 -> 4
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  19 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  18 <- 19
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  19 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,
  { b_lp ' (19) , b_lp ' (18) , b_lp ' (17) , b_lp ' (16)     }, // x =  0
  { b_lp ' (0) , b_lp ' (7) , b_lp ' (8) , b_lp ' (15)     }, // x =  1
  { b_lp ' (1) , b_lp ' (6) , b_lp ' (9) , b_lp ' (14)     }, // x =  2
  { b_lp ' (2) , b_lp ' (5) , b_lp ' (10) , b_lp ' (13)     }, // x =  3
  { b_lp ' (3) , b_lp ' (4) , b_lp ' (11) , b_lp ' (12)     } // x =  4
 };
end
if (x_max_p == 5  && y_max_p == 6 )
begin
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 4 ][ 5 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 4 ][ 5 ]; //  20 -> 21
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 3 ][ 5 ]; //  20 <- 21
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 3 ][ 5 ]; //  21 -> 22
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 2 ][ 5 ]; //  21 <- 22
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  22 <- 23
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 1 ][ 5 ]; //  23 -> 24
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 0 ][ 5 ]; //  23 <- 24
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 5 ]; //  24 -> 25
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 4 ][ 4 ]; //  18 <- 19
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 4 ][ 4 ]; //  19 -> 20
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 3 ][ 4 ]; //  17 <- 18
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 3 ][ 4 ]; //  18 -> 19
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 2 ][ 4 ]; //  16 <- 17
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 2 ][ 4 ]; //  17 -> 18
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 4 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 1 ][ 4 ]; //  16 -> 17
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 4 ]; //  24 <- 25
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 4 ]; //  25 -> 26
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  11 <- 12
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 4 ][ 3 ]; //  12 -> 13
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 3 ][ 3 ]; //  13 -> 14
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 2 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  14 <- 15
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 3 ]; //  15 -> 16
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 3 ]; //  25 <- 26
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  26 -> 27
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 4 ][ 2 ]; //  10 <- 11
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  11 -> 12
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 3 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  26 <- 27
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  27 -> 28
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 4 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  27 <- 28
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 4 ][ 0 ]; //  3 -> 4
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  29 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  28 <- 29
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  29 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,
  { b_lp ' (29) , b_lp ' (28) , b_lp ' (27) , b_lp ' (26) , b_lp ' (25) , b_lp ' (24)     }, // x =  0
  { b_lp ' (0) , b_lp ' (7) , b_lp ' (8) , b_lp ' (15) , b_lp ' (16) , b_lp ' (23)     }, // x =  1
  { b_lp ' (1) , b_lp ' (6) , b_lp ' (9) , b_lp ' (14) , b_lp ' (17) , b_lp ' (22)     }, // x =  2
  { b_lp ' (2) , b_lp ' (5) , b_lp ' (10) , b_lp ' (13) , b_lp ' (18) , b_lp ' (21)     }, // x =  3
  { b_lp ' (3) , b_lp ' (4) , b_lp ' (11) , b_lp ' (12) , b_lp ' (19) , b_lp ' (20)     } // x =  4
 };
end
if (x_max_p == 5  && y_max_p == 8 )
begin
assign back_data_in_o[ 4 ][ 6 ] = back_data_out_i[ 4 ][ 7 ]; //  27 <- 28
assign fwd_data_in_o [ 3 ][ 7 ] = fwd_data_out_i [ 4 ][ 7 ]; //  28 -> 29
assign back_data_in_o[ 4 ][ 7 ] = back_data_out_i[ 3 ][ 7 ]; //  28 <- 29
assign fwd_data_in_o [ 2 ][ 7 ] = fwd_data_out_i [ 3 ][ 7 ]; //  29 -> 30
assign back_data_in_o[ 3 ][ 7 ] = back_data_out_i[ 2 ][ 7 ]; //  29 <- 30
assign fwd_data_in_o [ 1 ][ 7 ] = fwd_data_out_i [ 2 ][ 7 ]; //  30 -> 31
assign back_data_in_o[ 2 ][ 7 ] = back_data_out_i[ 1 ][ 7 ]; //  30 <- 31
assign fwd_data_in_o [ 0 ][ 7 ] = fwd_data_out_i [ 1 ][ 7 ]; //  31 -> 32
assign back_data_in_o[ 1 ][ 7 ] = back_data_out_i[ 0 ][ 7 ]; //  31 <- 32
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 7 ]; //  32 -> 33
assign back_data_in_o[ 3 ][ 6 ] = back_data_out_i[ 4 ][ 6 ]; //  26 <- 27
assign fwd_data_in_o [ 4 ][ 7 ] = fwd_data_out_i [ 4 ][ 6 ]; //  27 -> 28
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 3 ][ 6 ]; //  25 <- 26
assign fwd_data_in_o [ 4 ][ 6 ] = fwd_data_out_i [ 3 ][ 6 ]; //  26 -> 27
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 2 ][ 6 ]; //  24 <- 25
assign fwd_data_in_o [ 3 ][ 6 ] = fwd_data_out_i [ 2 ][ 6 ]; //  25 -> 26
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 6 ]; //  23 <- 24
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 1 ][ 6 ]; //  24 -> 25
assign back_data_in_o[ 0 ][ 7 ] = back_data_out_i[ 0 ][ 6 ]; //  32 <- 33
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 6 ]; //  33 -> 34
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 4 ][ 5 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 4 ][ 5 ]; //  20 -> 21
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 3 ][ 5 ]; //  20 <- 21
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 3 ][ 5 ]; //  21 -> 22
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 2 ][ 5 ]; //  21 <- 22
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  22 <- 23
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 1 ][ 5 ]; //  23 -> 24
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 0 ][ 5 ]; //  33 <- 34
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 5 ]; //  34 -> 35
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 4 ][ 4 ]; //  18 <- 19
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 4 ][ 4 ]; //  19 -> 20
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 3 ][ 4 ]; //  17 <- 18
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 3 ][ 4 ]; //  18 -> 19
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 2 ][ 4 ]; //  16 <- 17
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 2 ][ 4 ]; //  17 -> 18
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 4 ]; //  15 <- 16
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 1 ][ 4 ]; //  16 -> 17
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 4 ]; //  34 <- 35
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 4 ]; //  35 -> 36
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 4 ][ 3 ]; //  11 <- 12
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 4 ][ 3 ]; //  12 -> 13
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  12 <- 13
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 3 ][ 3 ]; //  13 -> 14
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 2 ][ 3 ]; //  13 <- 14
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  14 -> 15
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  14 <- 15
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 3 ]; //  15 -> 16
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 3 ]; //  35 <- 36
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  36 -> 37
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 4 ][ 2 ]; //  10 <- 11
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 4 ][ 2 ]; //  11 -> 12
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  9 <- 10
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 3 ][ 2 ]; //  10 -> 11
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  8 <- 9
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  9 -> 10
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  7 <- 8
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  8 -> 9
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  36 <- 37
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  37 -> 38
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 4 ][ 1 ]; //  3 <- 4
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  4 -> 5
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  4 <- 5
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  5 -> 6
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  37 <- 38
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  38 -> 39
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 4 ][ 0 ]; //  3 -> 4
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  39 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  38 <- 39
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  39 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,  7,
  { b_lp ' (39) , b_lp ' (38) , b_lp ' (37) , b_lp ' (36) , b_lp ' (35) , b_lp ' (34) , b_lp ' (33) , b_lp ' (32)     }, // x =  0
  { b_lp ' (0) , b_lp ' (7) , b_lp ' (8) , b_lp ' (15) , b_lp ' (16) , b_lp ' (23) , b_lp ' (24) , b_lp ' (31)     }, // x =  1
  { b_lp ' (1) , b_lp ' (6) , b_lp ' (9) , b_lp ' (14) , b_lp ' (17) , b_lp ' (22) , b_lp ' (25) , b_lp ' (30)     }, // x =  2
  { b_lp ' (2) , b_lp ' (5) , b_lp ' (10) , b_lp ' (13) , b_lp ' (18) , b_lp ' (21) , b_lp ' (26) , b_lp ' (29)     }, // x =  3
  { b_lp ' (3) , b_lp ' (4) , b_lp ' (11) , b_lp ' (12) , b_lp ' (19) , b_lp ' (20) , b_lp ' (27) , b_lp ' (28)     } // x =  4
 };
end
if (x_max_p == 7  && y_max_p == 2 )
begin
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 6 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 6 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 5 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  9 -> 10
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 1 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 0 ][ 1 ]; //  11 <- 12
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  12 -> 13
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  4 <- 5
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 6 ][ 0 ]; //  5 -> 6
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  3 <- 4
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  4 -> 5
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  3 -> 4
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  13 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  12 <- 13
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  13 -> 0
 assign id_o =
 {
// y =  0,  1,
  { b_lp ' (13) , b_lp ' (12)     }, // x =  0
  { b_lp ' (0) , b_lp ' (11)     }, // x =  1
  { b_lp ' (1) , b_lp ' (10)     }, // x =  2
  { b_lp ' (2) , b_lp ' (9)     }, // x =  3
  { b_lp ' (3) , b_lp ' (8)     }, // x =  4
  { b_lp ' (4) , b_lp ' (7)     }, // x =  5
  { b_lp ' (5) , b_lp ' (6)     } // x =  6
 };
end
if (x_max_p == 7  && y_max_p == 4 )
begin
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 6 ][ 3 ]; //  17 <- 18
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 6 ][ 3 ]; //  18 -> 19
assign back_data_in_o[ 6 ][ 3 ] = back_data_out_i[ 5 ][ 3 ]; //  18 <- 19
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 5 ][ 3 ]; //  19 -> 20
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 4 ][ 3 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 4 ][ 3 ]; //  20 -> 21
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 3 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 2 ][ 3 ]; //  21 <- 22
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  22 <- 23
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 1 ][ 3 ]; //  23 -> 24
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 0 ][ 3 ]; //  23 <- 24
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  24 -> 25
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 6 ][ 2 ]; //  16 <- 17
assign fwd_data_in_o [ 6 ][ 3 ] = fwd_data_out_i [ 6 ][ 2 ]; //  17 -> 18
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 5 ][ 2 ]; //  15 <- 16
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 5 ][ 2 ]; //  16 -> 17
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 4 ][ 2 ]; //  14 <- 15
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 4 ][ 2 ]; //  15 -> 16
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  13 <- 14
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 3 ][ 2 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  12 -> 13
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  24 <- 25
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  25 -> 26
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 6 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 6 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 5 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  9 -> 10
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  25 <- 26
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  26 -> 27
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  4 <- 5
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 6 ][ 0 ]; //  5 -> 6
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  3 <- 4
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  4 -> 5
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  3 -> 4
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  27 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  26 <- 27
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  27 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,
  { b_lp ' (27) , b_lp ' (26) , b_lp ' (25) , b_lp ' (24)     }, // x =  0
  { b_lp ' (0) , b_lp ' (11) , b_lp ' (12) , b_lp ' (23)     }, // x =  1
  { b_lp ' (1) , b_lp ' (10) , b_lp ' (13) , b_lp ' (22)     }, // x =  2
  { b_lp ' (2) , b_lp ' (9) , b_lp ' (14) , b_lp ' (21)     }, // x =  3
  { b_lp ' (3) , b_lp ' (8) , b_lp ' (15) , b_lp ' (20)     }, // x =  4
  { b_lp ' (4) , b_lp ' (7) , b_lp ' (16) , b_lp ' (19)     }, // x =  5
  { b_lp ' (5) , b_lp ' (6) , b_lp ' (17) , b_lp ' (18)     } // x =  6
 };
end
if (x_max_p == 7  && y_max_p == 6 )
begin
assign back_data_in_o[ 6 ][ 4 ] = back_data_out_i[ 6 ][ 5 ]; //  29 <- 30
assign fwd_data_in_o [ 5 ][ 5 ] = fwd_data_out_i [ 6 ][ 5 ]; //  30 -> 31
assign back_data_in_o[ 6 ][ 5 ] = back_data_out_i[ 5 ][ 5 ]; //  30 <- 31
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 5 ][ 5 ]; //  31 -> 32
assign back_data_in_o[ 5 ][ 5 ] = back_data_out_i[ 4 ][ 5 ]; //  31 <- 32
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 4 ][ 5 ]; //  32 -> 33
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 3 ][ 5 ]; //  32 <- 33
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 3 ][ 5 ]; //  33 -> 34
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 2 ][ 5 ]; //  33 <- 34
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  34 -> 35
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  34 <- 35
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 1 ][ 5 ]; //  35 -> 36
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 0 ][ 5 ]; //  35 <- 36
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 5 ]; //  36 -> 37
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 6 ][ 4 ]; //  28 <- 29
assign fwd_data_in_o [ 6 ][ 5 ] = fwd_data_out_i [ 6 ][ 4 ]; //  29 -> 30
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 5 ][ 4 ]; //  27 <- 28
assign fwd_data_in_o [ 6 ][ 4 ] = fwd_data_out_i [ 5 ][ 4 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 4 ][ 4 ]; //  26 <- 27
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 4 ][ 4 ]; //  27 -> 28
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 3 ][ 4 ]; //  25 <- 26
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 3 ][ 4 ]; //  26 -> 27
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 2 ][ 4 ]; //  24 <- 25
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 2 ][ 4 ]; //  25 -> 26
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 4 ]; //  23 <- 24
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 1 ][ 4 ]; //  24 -> 25
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 4 ]; //  36 <- 37
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 4 ]; //  37 -> 38
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 6 ][ 3 ]; //  17 <- 18
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 6 ][ 3 ]; //  18 -> 19
assign back_data_in_o[ 6 ][ 3 ] = back_data_out_i[ 5 ][ 3 ]; //  18 <- 19
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 5 ][ 3 ]; //  19 -> 20
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 4 ][ 3 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 4 ][ 3 ]; //  20 -> 21
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 3 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 2 ][ 3 ]; //  21 <- 22
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  22 <- 23
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 3 ]; //  23 -> 24
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 3 ]; //  37 <- 38
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  38 -> 39
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 6 ][ 2 ]; //  16 <- 17
assign fwd_data_in_o [ 6 ][ 3 ] = fwd_data_out_i [ 6 ][ 2 ]; //  17 -> 18
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 5 ][ 2 ]; //  15 <- 16
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 5 ][ 2 ]; //  16 -> 17
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 4 ][ 2 ]; //  14 <- 15
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 4 ][ 2 ]; //  15 -> 16
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  13 <- 14
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 3 ][ 2 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  12 -> 13
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  38 <- 39
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  39 -> 40
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 6 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 6 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 5 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  9 -> 10
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  39 <- 40
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  40 -> 41
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  4 <- 5
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 6 ][ 0 ]; //  5 -> 6
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  3 <- 4
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  4 -> 5
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  3 -> 4
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  41 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  40 <- 41
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  41 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,
  { b_lp ' (41) , b_lp ' (40) , b_lp ' (39) , b_lp ' (38) , b_lp ' (37) , b_lp ' (36)     }, // x =  0
  { b_lp ' (0) , b_lp ' (11) , b_lp ' (12) , b_lp ' (23) , b_lp ' (24) , b_lp ' (35)     }, // x =  1
  { b_lp ' (1) , b_lp ' (10) , b_lp ' (13) , b_lp ' (22) , b_lp ' (25) , b_lp ' (34)     }, // x =  2
  { b_lp ' (2) , b_lp ' (9) , b_lp ' (14) , b_lp ' (21) , b_lp ' (26) , b_lp ' (33)     }, // x =  3
  { b_lp ' (3) , b_lp ' (8) , b_lp ' (15) , b_lp ' (20) , b_lp ' (27) , b_lp ' (32)     }, // x =  4
  { b_lp ' (4) , b_lp ' (7) , b_lp ' (16) , b_lp ' (19) , b_lp ' (28) , b_lp ' (31)     }, // x =  5
  { b_lp ' (5) , b_lp ' (6) , b_lp ' (17) , b_lp ' (18) , b_lp ' (29) , b_lp ' (30)     } // x =  6
 };
end
if (x_max_p == 7  && y_max_p == 8 )
begin
assign back_data_in_o[ 6 ][ 6 ] = back_data_out_i[ 6 ][ 7 ]; //  41 <- 42
assign fwd_data_in_o [ 5 ][ 7 ] = fwd_data_out_i [ 6 ][ 7 ]; //  42 -> 43
assign back_data_in_o[ 6 ][ 7 ] = back_data_out_i[ 5 ][ 7 ]; //  42 <- 43
assign fwd_data_in_o [ 4 ][ 7 ] = fwd_data_out_i [ 5 ][ 7 ]; //  43 -> 44
assign back_data_in_o[ 5 ][ 7 ] = back_data_out_i[ 4 ][ 7 ]; //  43 <- 44
assign fwd_data_in_o [ 3 ][ 7 ] = fwd_data_out_i [ 4 ][ 7 ]; //  44 -> 45
assign back_data_in_o[ 4 ][ 7 ] = back_data_out_i[ 3 ][ 7 ]; //  44 <- 45
assign fwd_data_in_o [ 2 ][ 7 ] = fwd_data_out_i [ 3 ][ 7 ]; //  45 -> 46
assign back_data_in_o[ 3 ][ 7 ] = back_data_out_i[ 2 ][ 7 ]; //  45 <- 46
assign fwd_data_in_o [ 1 ][ 7 ] = fwd_data_out_i [ 2 ][ 7 ]; //  46 -> 47
assign back_data_in_o[ 2 ][ 7 ] = back_data_out_i[ 1 ][ 7 ]; //  46 <- 47
assign fwd_data_in_o [ 0 ][ 7 ] = fwd_data_out_i [ 1 ][ 7 ]; //  47 -> 48
assign back_data_in_o[ 1 ][ 7 ] = back_data_out_i[ 0 ][ 7 ]; //  47 <- 48
assign fwd_data_in_o [ 0 ][ 6 ] = fwd_data_out_i [ 0 ][ 7 ]; //  48 -> 49
assign back_data_in_o[ 5 ][ 6 ] = back_data_out_i[ 6 ][ 6 ]; //  40 <- 41
assign fwd_data_in_o [ 6 ][ 7 ] = fwd_data_out_i [ 6 ][ 6 ]; //  41 -> 42
assign back_data_in_o[ 4 ][ 6 ] = back_data_out_i[ 5 ][ 6 ]; //  39 <- 40
assign fwd_data_in_o [ 6 ][ 6 ] = fwd_data_out_i [ 5 ][ 6 ]; //  40 -> 41
assign back_data_in_o[ 3 ][ 6 ] = back_data_out_i[ 4 ][ 6 ]; //  38 <- 39
assign fwd_data_in_o [ 5 ][ 6 ] = fwd_data_out_i [ 4 ][ 6 ]; //  39 -> 40
assign back_data_in_o[ 2 ][ 6 ] = back_data_out_i[ 3 ][ 6 ]; //  37 <- 38
assign fwd_data_in_o [ 4 ][ 6 ] = fwd_data_out_i [ 3 ][ 6 ]; //  38 -> 39
assign back_data_in_o[ 1 ][ 6 ] = back_data_out_i[ 2 ][ 6 ]; //  36 <- 37
assign fwd_data_in_o [ 3 ][ 6 ] = fwd_data_out_i [ 2 ][ 6 ]; //  37 -> 38
assign back_data_in_o[ 1 ][ 5 ] = back_data_out_i[ 1 ][ 6 ]; //  35 <- 36
assign fwd_data_in_o [ 2 ][ 6 ] = fwd_data_out_i [ 1 ][ 6 ]; //  36 -> 37
assign back_data_in_o[ 0 ][ 7 ] = back_data_out_i[ 0 ][ 6 ]; //  48 <- 49
assign fwd_data_in_o [ 0 ][ 5 ] = fwd_data_out_i [ 0 ][ 6 ]; //  49 -> 50
assign back_data_in_o[ 6 ][ 4 ] = back_data_out_i[ 6 ][ 5 ]; //  29 <- 30
assign fwd_data_in_o [ 5 ][ 5 ] = fwd_data_out_i [ 6 ][ 5 ]; //  30 -> 31
assign back_data_in_o[ 6 ][ 5 ] = back_data_out_i[ 5 ][ 5 ]; //  30 <- 31
assign fwd_data_in_o [ 4 ][ 5 ] = fwd_data_out_i [ 5 ][ 5 ]; //  31 -> 32
assign back_data_in_o[ 5 ][ 5 ] = back_data_out_i[ 4 ][ 5 ]; //  31 <- 32
assign fwd_data_in_o [ 3 ][ 5 ] = fwd_data_out_i [ 4 ][ 5 ]; //  32 -> 33
assign back_data_in_o[ 4 ][ 5 ] = back_data_out_i[ 3 ][ 5 ]; //  32 <- 33
assign fwd_data_in_o [ 2 ][ 5 ] = fwd_data_out_i [ 3 ][ 5 ]; //  33 -> 34
assign back_data_in_o[ 3 ][ 5 ] = back_data_out_i[ 2 ][ 5 ]; //  33 <- 34
assign fwd_data_in_o [ 1 ][ 5 ] = fwd_data_out_i [ 2 ][ 5 ]; //  34 -> 35
assign back_data_in_o[ 2 ][ 5 ] = back_data_out_i[ 1 ][ 5 ]; //  34 <- 35
assign fwd_data_in_o [ 1 ][ 6 ] = fwd_data_out_i [ 1 ][ 5 ]; //  35 -> 36
assign back_data_in_o[ 0 ][ 6 ] = back_data_out_i[ 0 ][ 5 ]; //  49 <- 50
assign fwd_data_in_o [ 0 ][ 4 ] = fwd_data_out_i [ 0 ][ 5 ]; //  50 -> 51
assign back_data_in_o[ 5 ][ 4 ] = back_data_out_i[ 6 ][ 4 ]; //  28 <- 29
assign fwd_data_in_o [ 6 ][ 5 ] = fwd_data_out_i [ 6 ][ 4 ]; //  29 -> 30
assign back_data_in_o[ 4 ][ 4 ] = back_data_out_i[ 5 ][ 4 ]; //  27 <- 28
assign fwd_data_in_o [ 6 ][ 4 ] = fwd_data_out_i [ 5 ][ 4 ]; //  28 -> 29
assign back_data_in_o[ 3 ][ 4 ] = back_data_out_i[ 4 ][ 4 ]; //  26 <- 27
assign fwd_data_in_o [ 5 ][ 4 ] = fwd_data_out_i [ 4 ][ 4 ]; //  27 -> 28
assign back_data_in_o[ 2 ][ 4 ] = back_data_out_i[ 3 ][ 4 ]; //  25 <- 26
assign fwd_data_in_o [ 4 ][ 4 ] = fwd_data_out_i [ 3 ][ 4 ]; //  26 -> 27
assign back_data_in_o[ 1 ][ 4 ] = back_data_out_i[ 2 ][ 4 ]; //  24 <- 25
assign fwd_data_in_o [ 3 ][ 4 ] = fwd_data_out_i [ 2 ][ 4 ]; //  25 -> 26
assign back_data_in_o[ 1 ][ 3 ] = back_data_out_i[ 1 ][ 4 ]; //  23 <- 24
assign fwd_data_in_o [ 2 ][ 4 ] = fwd_data_out_i [ 1 ][ 4 ]; //  24 -> 25
assign back_data_in_o[ 0 ][ 5 ] = back_data_out_i[ 0 ][ 4 ]; //  50 <- 51
assign fwd_data_in_o [ 0 ][ 3 ] = fwd_data_out_i [ 0 ][ 4 ]; //  51 -> 52
assign back_data_in_o[ 6 ][ 2 ] = back_data_out_i[ 6 ][ 3 ]; //  17 <- 18
assign fwd_data_in_o [ 5 ][ 3 ] = fwd_data_out_i [ 6 ][ 3 ]; //  18 -> 19
assign back_data_in_o[ 6 ][ 3 ] = back_data_out_i[ 5 ][ 3 ]; //  18 <- 19
assign fwd_data_in_o [ 4 ][ 3 ] = fwd_data_out_i [ 5 ][ 3 ]; //  19 -> 20
assign back_data_in_o[ 5 ][ 3 ] = back_data_out_i[ 4 ][ 3 ]; //  19 <- 20
assign fwd_data_in_o [ 3 ][ 3 ] = fwd_data_out_i [ 4 ][ 3 ]; //  20 -> 21
assign back_data_in_o[ 4 ][ 3 ] = back_data_out_i[ 3 ][ 3 ]; //  20 <- 21
assign fwd_data_in_o [ 2 ][ 3 ] = fwd_data_out_i [ 3 ][ 3 ]; //  21 -> 22
assign back_data_in_o[ 3 ][ 3 ] = back_data_out_i[ 2 ][ 3 ]; //  21 <- 22
assign fwd_data_in_o [ 1 ][ 3 ] = fwd_data_out_i [ 2 ][ 3 ]; //  22 -> 23
assign back_data_in_o[ 2 ][ 3 ] = back_data_out_i[ 1 ][ 3 ]; //  22 <- 23
assign fwd_data_in_o [ 1 ][ 4 ] = fwd_data_out_i [ 1 ][ 3 ]; //  23 -> 24
assign back_data_in_o[ 0 ][ 4 ] = back_data_out_i[ 0 ][ 3 ]; //  51 <- 52
assign fwd_data_in_o [ 0 ][ 2 ] = fwd_data_out_i [ 0 ][ 3 ]; //  52 -> 53
assign back_data_in_o[ 5 ][ 2 ] = back_data_out_i[ 6 ][ 2 ]; //  16 <- 17
assign fwd_data_in_o [ 6 ][ 3 ] = fwd_data_out_i [ 6 ][ 2 ]; //  17 -> 18
assign back_data_in_o[ 4 ][ 2 ] = back_data_out_i[ 5 ][ 2 ]; //  15 <- 16
assign fwd_data_in_o [ 6 ][ 2 ] = fwd_data_out_i [ 5 ][ 2 ]; //  16 -> 17
assign back_data_in_o[ 3 ][ 2 ] = back_data_out_i[ 4 ][ 2 ]; //  14 <- 15
assign fwd_data_in_o [ 5 ][ 2 ] = fwd_data_out_i [ 4 ][ 2 ]; //  15 -> 16
assign back_data_in_o[ 2 ][ 2 ] = back_data_out_i[ 3 ][ 2 ]; //  13 <- 14
assign fwd_data_in_o [ 4 ][ 2 ] = fwd_data_out_i [ 3 ][ 2 ]; //  14 -> 15
assign back_data_in_o[ 1 ][ 2 ] = back_data_out_i[ 2 ][ 2 ]; //  12 <- 13
assign fwd_data_in_o [ 3 ][ 2 ] = fwd_data_out_i [ 2 ][ 2 ]; //  13 -> 14
assign back_data_in_o[ 1 ][ 1 ] = back_data_out_i[ 1 ][ 2 ]; //  11 <- 12
assign fwd_data_in_o [ 2 ][ 2 ] = fwd_data_out_i [ 1 ][ 2 ]; //  12 -> 13
assign back_data_in_o[ 0 ][ 3 ] = back_data_out_i[ 0 ][ 2 ]; //  52 <- 53
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 2 ]; //  53 -> 54
assign back_data_in_o[ 6 ][ 0 ] = back_data_out_i[ 6 ][ 1 ]; //  5 <- 6
assign fwd_data_in_o [ 5 ][ 1 ] = fwd_data_out_i [ 6 ][ 1 ]; //  6 -> 7
assign back_data_in_o[ 6 ][ 1 ] = back_data_out_i[ 5 ][ 1 ]; //  6 <- 7
assign fwd_data_in_o [ 4 ][ 1 ] = fwd_data_out_i [ 5 ][ 1 ]; //  7 -> 8
assign back_data_in_o[ 5 ][ 1 ] = back_data_out_i[ 4 ][ 1 ]; //  7 <- 8
assign fwd_data_in_o [ 3 ][ 1 ] = fwd_data_out_i [ 4 ][ 1 ]; //  8 -> 9
assign back_data_in_o[ 4 ][ 1 ] = back_data_out_i[ 3 ][ 1 ]; //  8 <- 9
assign fwd_data_in_o [ 2 ][ 1 ] = fwd_data_out_i [ 3 ][ 1 ]; //  9 -> 10
assign back_data_in_o[ 3 ][ 1 ] = back_data_out_i[ 2 ][ 1 ]; //  9 <- 10
assign fwd_data_in_o [ 1 ][ 1 ] = fwd_data_out_i [ 2 ][ 1 ]; //  10 -> 11
assign back_data_in_o[ 2 ][ 1 ] = back_data_out_i[ 1 ][ 1 ]; //  10 <- 11
assign fwd_data_in_o [ 1 ][ 2 ] = fwd_data_out_i [ 1 ][ 1 ]; //  11 -> 12
assign back_data_in_o[ 0 ][ 2 ] = back_data_out_i[ 0 ][ 1 ]; //  53 <- 54
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  54 -> 55
assign back_data_in_o[ 5 ][ 0 ] = back_data_out_i[ 6 ][ 0 ]; //  4 <- 5
assign fwd_data_in_o [ 6 ][ 1 ] = fwd_data_out_i [ 6 ][ 0 ]; //  5 -> 6
assign back_data_in_o[ 4 ][ 0 ] = back_data_out_i[ 5 ][ 0 ]; //  3 <- 4
assign fwd_data_in_o [ 6 ][ 0 ] = fwd_data_out_i [ 5 ][ 0 ]; //  4 -> 5
assign back_data_in_o[ 3 ][ 0 ] = back_data_out_i[ 4 ][ 0 ]; //  2 <- 3
assign fwd_data_in_o [ 5 ][ 0 ] = fwd_data_out_i [ 4 ][ 0 ]; //  3 -> 4
assign back_data_in_o[ 2 ][ 0 ] = back_data_out_i[ 3 ][ 0 ]; //  1 <- 2
assign fwd_data_in_o [ 4 ][ 0 ] = fwd_data_out_i [ 3 ][ 0 ]; //  2 -> 3
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 2 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 3 ][ 0 ] = fwd_data_out_i [ 2 ][ 0 ]; //  1 -> 2
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  55 <- 0
assign fwd_data_in_o [ 2 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  0 -> 1
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  54 <- 55
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  55 -> 0
 assign id_o =
 {
// y =  0,  1,  2,  3,  4,  5,  6,  7,
  { b_lp ' (55) , b_lp ' (54) , b_lp ' (53) , b_lp ' (52) , b_lp ' (51) , b_lp ' (50) , b_lp ' (49) , b_lp ' (48)     }, // x =  0
  { b_lp ' (0) , b_lp ' (11) , b_lp ' (12) , b_lp ' (23) , b_lp ' (24) , b_lp ' (35) , b_lp ' (36) , b_lp ' (47)     }, // x =  1
  { b_lp ' (1) , b_lp ' (10) , b_lp ' (13) , b_lp ' (22) , b_lp ' (25) , b_lp ' (34) , b_lp ' (37) , b_lp ' (46)     }, // x =  2
  { b_lp ' (2) , b_lp ' (9) , b_lp ' (14) , b_lp ' (21) , b_lp ' (26) , b_lp ' (33) , b_lp ' (38) , b_lp ' (45)     }, // x =  3
  { b_lp ' (3) , b_lp ' (8) , b_lp ' (15) , b_lp ' (20) , b_lp ' (27) , b_lp ' (32) , b_lp ' (39) , b_lp ' (44)     }, // x =  4
  { b_lp ' (4) , b_lp ' (7) , b_lp ' (16) , b_lp ' (19) , b_lp ' (28) , b_lp ' (31) , b_lp ' (40) , b_lp ' (43)     }, // x =  5
  { b_lp ' (5) , b_lp ' (6) , b_lp ' (17) , b_lp ' (18) , b_lp ' (29) , b_lp ' (30) , b_lp ' (41) , b_lp ' (42)     } // x =  6
 };
end
if (x_max_p == 1  && y_max_p == 2 )
begin
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 0 ][ 1 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 0 ][ 1 ]; //  1 -> 0
assign back_data_in_o[ 0 ][ 1 ] = back_data_out_i[ 0 ][ 0 ]; //  1 <- 0
assign fwd_data_in_o [ 0 ][ 1 ] = fwd_data_out_i [ 0 ][ 0 ]; //  0 -> 1
 assign id_o =
 {
// y =  0,  1,
  { b_lp ' (0) , b_lp ' (1)     } // x =  0
 };
end
if (x_max_p == 2  && y_max_p == 1 )
begin
assign back_data_in_o[ 0 ][ 0 ] = back_data_out_i[ 1 ][ 0 ]; //  0 <- 1
assign fwd_data_in_o [ 0 ][ 0 ] = fwd_data_out_i [ 1 ][ 0 ]; //  1 -> 0
assign back_data_in_o[ 1 ][ 0 ] = back_data_out_i[ 0 ][ 0 ]; //  1 <- 0
assign fwd_data_in_o [ 1 ][ 0 ] = fwd_data_out_i [ 0 ][ 0 ]; //  0 -> 1
 assign id_o =
 {
// y =  0,
  { b_lp ' (0)     }, // x =  0
  { b_lp ' (1)     } // x =  1
 };
end
initial assert ((x_max_p <= 8) && (y_max_p <= 8)) else begin $error("%m x_max_p %d or y_max_p %d too large; rerun generator with larger size than %d/%d",x_max_p,y_max_p,8,8); $finish(); end
endmodule