module xsv_fpga_top (
	// Global signals
	clk, rstn, /*tx_clk, rx_clk,*/
	// Flash chip
	flash_rstn, flash_cen, flash_oen, flash_wen,
	flash_rdy, flash_d, flash_a,
	// SRAM right bank
	sram_r_cen, sram_r_oen, sram_r0_wen,
	sram_r1_wen, sram_r_d, sram_r_a,
	// SRAM left bank
	sram_l_cen, sram_l_oen, sram_l0_wen,
	sram_l1_wen, sram_l_d, sram_l_a,
	`ifdef SPOOFER
	clk_count,spoof_out,trigger,
	`endif
/*
`ifdef APP_VGA_RAMDAC
	// VGA RAMDAC
	ramdac_pixclk, ramdac_hsyncn, ramdac_vsync, ramdac_blank,
	ramdac_p, ramdac_rdn, ramdac_wrn, ramdac_rs, ramdac_d,
`else
	// VGA Direct
	vga_blank, vga_pclk, vga_hsyncn, vga_vsyncn,
	vga_r, vga_g, vga_b,
`endif
	// Stereo Codec
	codec_mclk, codec_lrclk, codec_sclk,
	codec_sdin, codec_sdout,
*/
/*
	// Ethernet
	eth_col, eth_crs, eth_trste, eth_tx_clk,
	eth_tx_en, eth_tx_er, eth_txd, eth_rx_clk,
	eth_rx_dv, eth_rx_er, eth_rxd, eth_fds_mdint,
	eth_mdc, eth_mdio,
*/
	// Switches
	sw,
/*
	// PS/2 keyboard
	ps2_clk, ps2_data,
*/
	// CPLD
	tdmfrm, tdmrx, tdmtx
);
// I/O Ports
// Global
input			clk;
input			rstn;
/*
input    tx_clk;
input    rx_clk;
*/
// Flash
output 			flash_rstn;
output 			flash_cen;
output 			flash_oen;
output 			flash_wen;
input 			flash_rdy;
inout	[7:0]		flash_d;
inout	[20:0]		flash_a;
// SRAM Right
output			sram_r_cen;
output			sram_r1_wen;
output			sram_r0_wen;
output			sram_r_oen;
output	[18:0]		sram_r_a;
inout	[15:0]		sram_r_d;
// SRAM Left
output			sram_l_cen;
output			sram_l0_wen;
output			sram_l1_wen;
output			sram_l_oen;
output	[18:0]		sram_l_a;
inout	[15:0]		sram_l_d;
`ifdef SPOOFER
input	[31:0]		clk_count;
output	[31:0]		spoof_out;
output			trigger;
`endif
/*
`ifdef APP_VGA_RAMDAC
// VGA RAMDAC
output			ramdac_pixclk;
output			ramdac_hsyncn;
output			ramdac_vsync;
output			ramdac_blank;
output	[7:0]		ramdac_p;
output			ramdac_rdn;
output			ramdac_wrn;
output	[2:0]		ramdac_rs;
inout	[7:0]		ramdac_d;
`else
// VGA Direct
output			vga_pclk;
output			vga_blank;
output			vga_hsyncn;
output			vga_vsyncn;
output	[3:0]		vga_r;
output	[3:0]		vga_g;
output	[3:0]		vga_b;
`endif
// Stereo Codec
output			codec_mclk;
output			codec_lrclk;
output			codec_sclk;
output			codec_sdin;
input			codec_sdout;
*/
/*
// Ethernet
output			eth_tx_er;
input			eth_tx_clk;
output			eth_tx_en;
output	[3:0]		eth_txd;
input			eth_rx_er;
input			eth_rx_clk;
input			eth_rx_dv;
input	[3:0]		eth_rxd;
input			eth_col;
input			eth_crs;
output			eth_trste;
input			eth_fds_mdint;
inout			eth_mdio;
output			eth_mdc;
*/
// Switches
input	[2:1]		sw;
/*
// PS/2 keyboard
inout			ps2_clk;
inout			ps2_data;
*/
// CPLD TDM
input			tdmfrm;
input			tdmrx;
output			tdmtx;
// Internal wires
/*
// VGA core slave i/f wires
wire 	[31:0]		wb_vs_adr_i;
wire 	[31:0]		wb_vs_dat_i;
wire 	[31:0]		wb_vs_dat_o;
wire 	[3:0]		wb_vs_sel_i;
wire 			wb_vs_we_i;
wire 			wb_vs_stb_i;
wire 			wb_vs_cyc_i;
wire 			wb_vs_ack_o;
wire 			wb_vs_err_o;
// VGA core master i/f wires
wire 	[31:0]		wb_vm_adr_o;
wire 	[31:0] 		wb_vm_dat_i;
wire 	[3:0]		wb_vm_sel_o;
wire			wb_vm_we_o;
wire 			wb_vm_stb_o;
wire			wb_vm_cyc_o;
wire			wb_vm_cab_o;
wire			wb_vm_ack_i;
wire			wb_vm_err_i;
// VGA CRT wires
wire	[4:0]		vga_r_int;
wire	[5:0]		vga_g_int;
wire	[4:0]		vga_b_int;
wire			crt_hsync;
wire			crt_vsync;
*/
`ifdef SPOOFER
wire	[31:0]   	clk_count;
wire  	[31:0]		spoof_out;
wire			trigger;
`endif
// Debug core master i/f wires
wire 	[31:0]		wb_dm_adr_o;
wire 	[31:0] 		wb_dm_dat_i;
wire 	[31:0] 		wb_dm_dat_o;
wire 	[3:0]		wb_dm_sel_o;
wire			wb_dm_we_o;
wire 			wb_dm_stb_o;
wire			wb_dm_cyc_o;
wire			wb_dm_cab_o;
wire			wb_dm_ack_i;
wire			wb_dm_err_i;
// Debug <-> RISC wires
wire	[3:0]		dbg_lss;
wire	[1:0]		dbg_is;
wire	[10:0]		dbg_wp;
wire			dbg_bp;
wire	[31:0]		dbg_dat_dbg;
wire	[31:0]		dbg_dat_risc;
wire	[31:0]		dbg_adr;
wire			dbg_ewt;
wire			dbg_stall;
wire	[2:0]		dbg_op;
// RISC instruction master i/f wires
wire 	[31:0]		wb_rim_adr_o;
wire			wb_rim_cyc_o;
wire 	[31:0]		wb_rim_dat_i;
wire 	[31:0]		wb_rim_dat_o;
wire 	[3:0]		wb_rim_sel_o;
wire			wb_rim_ack_i;
wire			wb_rim_err_i;
wire			wb_rim_rty_i = 1'b0;
wire			wb_rim_we_o;
wire			wb_rim_stb_o;
wire			wb_rim_cab_o;
wire	[31:0]		wb_rif_adr;
reg			prefix_flash;
// RISC data master i/f wires
wire 	[31:0]		wb_rdm_adr_o;
wire			wb_rdm_cyc_o;
wire 	[31:0]		wb_rdm_dat_i;
wire 	[31:0]		wb_rdm_dat_o;
wire 	[3:0]		wb_rdm_sel_o;
wire			wb_rdm_ack_i;
wire			wb_rdm_err_i;
wire			wb_rdm_rty_i = 1'b0;
wire			wb_rdm_we_o;
wire			wb_rdm_stb_o;
wire			wb_rdm_cab_o;
wire			wb_rdm_ack;
// RISC misc
wire	[19:0]		pic_ints;
// SRAM controller slave i/f wires
wire 	[31:0]		wb_ss_dat_i;
wire 	[31:0]		wb_ss_dat_o;
wire 	[31:0]		wb_ss_adr_i;
wire 	[3:0]		wb_ss_sel_i;
wire			wb_ss_we_i;
wire			wb_ss_cyc_i;
wire			wb_ss_stb_i;
wire			wb_ss_ack_o;
wire			wb_ss_err_o;
// SRAM external wires
wire	[15:0]		sram_r_d_o;
wire	[15:0]		sram_l_d_o;
wire			sram_d_oe;
// Flash controller slave i/f wires
wire 	[31:0]		wb_fs_dat_i;
wire 	[31:0]		wb_fs_dat_o;
wire 	[31:0]		wb_fs_adr_i;
wire 	[3:0]		wb_fs_sel_i;
wire			wb_fs_we_i;
wire			wb_fs_cyc_i;
wire			wb_fs_stb_i;
wire			wb_fs_ack_o;
wire			wb_fs_err_o;
/*
// Audio core slave i/f wires
wire 	[31:0]		wb_as_dat_i;
wire 	[31:0]		wb_as_dat_o;
wire 	[31:0]		wb_as_adr_i;
wire 	[3:0]		wb_as_sel_i;
wire			wb_as_we_i;
wire			wb_as_cyc_i;
wire			wb_as_stb_i;
wire			wb_as_ack_o;
wire			wb_as_err_o;
// Audio core master i/f wires
wire 	[31:0]		wb_am_dat_o;
wire 	[31:0]		wb_am_dat_i;
wire 	[31:0]		wb_am_adr_o;
wire 	[3:0]		wb_am_sel_o;
wire			wb_am_we_o;
wire			wb_am_cyc_o;
wire			wb_am_stb_o;
wire			wb_am_cab_o;
wire			wb_am_ack_i;
wire			wb_am_err_i;
// PS/2 core slave i/f wires
wire 	[31:0]		wb_ps_dat_i;
wire 	[31:0]		wb_ps_dat_o;
wire 	[31:0]		wb_ps_adr_i;
wire 	[3:0]		wb_ps_sel_i;
wire			wb_ps_we_i;
wire			wb_ps_cyc_i;
wire			wb_ps_stb_i;
wire			wb_ps_ack_o;
wire			wb_ps_err_o;
// PS/2 external i/f wires
wire			ps2_clk_o;
wire			ps2_data_o;
wire			ps2_clk_oe;
wire			ps2_data_oe;
// Ethernet core master i/f wires
wire 	[31:0]		wb_em_adr_o;
wire 	[31:0] 		wb_em_dat_i;
wire 	[31:0] 		wb_em_dat_o;
wire 	[3:0]		wb_em_sel_o;
wire			wb_em_we_o;
wire 			wb_em_stb_o;
wire			wb_em_cyc_o;
wire			wb_em_cab_o;
wire			wb_em_ack_i;
wire			wb_em_err_i;
// Ethernet core slave i/f wires
wire	[31:0]		wb_es_dat_i;
wire	[31:0]		wb_es_dat_o;
wire	[31:0]		wb_es_adr_i;
wire	[3:0]		wb_es_sel_i;
wire			wb_es_we_i;
wire			wb_es_cyc_i;
wire			wb_es_stb_i;
wire			wb_es_ack_o;
wire			wb_es_err_o;
// Ethernet external i/f wires
wire			eth_mdo;
wire			eth_mdoe;
// UART16550 core slave i/f wires
wire	[31:0]		wb_us_dat_i;
wire	[31:0]		wb_us_dat_o;
wire	[31:0]		wb_us_adr_i;
wire	[3:0]		wb_us_sel_i;
wire			wb_us_we_i;
wire			wb_us_cyc_i;
wire			wb_us_stb_i;
wire			wb_us_ack_o;
wire			wb_us_err_o;
// HDLC core slave i/f wires
//wire	[31:0]		wb_hd_dat_i;
//wire	[31:0]		wb_hd_dat_o;
//wire	[31:0]		wb_hd_adr_i;
//wire	[3:0]		wb_hd_sel_i;
//wire			wb_hd_we_i;
//wire			wb_hd_cyc_i;
//wire			wb_hd_stb_i;
//wire			wb_hd_ack_o;
//wire			wb_hd_err_o;
//wire     tx_clk;
//wire     rx_clk;
// HDLC external i/f wires
//wire			hdlc_tx;
//wire			hdlc_rx;
//wire     Loopback;
// UART external i/f wires
//wire			uart_stx;
//wire			uart_srx;
*/
// JTAG wires
wire			jtag_tdi;
wire			jtag_tms;
wire			jtag_tck;
wire			jtag_trst;
wire			jtag_tdo;
// CPLD TDM wires
wire	[2:0]		tdm_out_unused;
reg  [2:0] wb_hd_adr_i_map;
// Reset debounce
reg			rst_r;
reg			wb_rst;
// Global clock
`ifdef OR1200_CLMODE_1TO2
reg			wb_clk;
`else
wire			wb_clk;
`endif
// Reset debounce
always @(posedge wb_clk or negedge rstn)
	if (~rstn)
		rst_r <= 1'b1;
	else
		rst_r <= #1 1'b0;
// Reset debounce
always @(posedge wb_clk)
	wb_rst <= #1 rst_r;
// This is purely for testing 1/2 WB clock
// This should never be used when implementing in
// an FPGA. It is used only for simulation regressions.
`ifdef OR1200_CLMODE_1TO2
initial wb_clk = 0;
always @(posedge clk)
	wb_clk = ~wb_clk;
`else
// Some Xilinx P&R tools need this
`ifdef TARGET_VIRTEX
IBUFG IBUFG1 (
	.O	( wb_clk ),
	.I	( clk )
);
`else
assign wb_clk = clk;
`endif
`endif // OR1200_CLMODE_1TO2
// SRAM tri-state data
assign sram_r_d = sram_d_oe ? sram_r_d_o : 16'hzzzz;
assign sram_l_d = sram_d_oe ? sram_l_d_o : 16'hzzzz;
// Ethernet tri-state
//assign eth_mdio = eth_mdoe ? eth_mdo : 1'bz;
//assign eth_trste = 1'b0;
// PS/2 Keyboard tri-state
//assign ps2_clk = ps2_clk_oe ? ps2_clk_o : 1'bz;
//assign ps2_data = ps2_data_oe ? ps2_data_o : 1'bz;
// Unused interrupts
/*assign pic_ints[`APP_INT_RES1] = 'b0;
assign pic_ints[`APP_INT_RES2] = 'b0;
assign pic_ints[`APP_INT_RES3] = 'b0;*/
assign pic_ints[19:0] = 20'b0;
// Unused WISHBONE signals
assign wb_hd_err_o = 1'b0;
assign wb_us_err_o = 1'b0;
assign wb_ps_err_o = 1'b0;
assign wb_em_cab_o = 1'b0;
assign wb_am_cab_o = 1'b0;
// RISC Instruction address for Flash
// Until first access to real Flash area,
// it is always prefixed with Flash area prefix.
// This way we have flash at base address 0x0
// during reset vector execution (boot). First
// access to real Flash area will automatically
// move SRAM to 0x0.
always @(posedge wb_clk or negedge rstn)
	if (!rstn)
		prefix_flash <= #1 1'b1;
	else if (wb_rim_cyc_o &&
		(wb_rim_adr_o[31:32-`APP_ADDR_DEC_W] == `APP_ADDR_FLASH))
		prefix_flash <= #1 1'b0;
assign wb_rif_adr = prefix_flash ? {`APP_ADDR_FLASH, wb_rim_adr_o[31-`APP_ADDR_DEC_W:0]}
			: wb_rim_adr_o;
assign wb_rdm_ack_i = (wb_rdm_adr_o[31:28] == `APP_ADDR_FAKEMC) &&
			wb_rdm_cyc_o && wb_rdm_stb_o ? 1'b1 : wb_rdm_ack;
// Instantiation of the VGA CRT controller
/*
ssvga_top ssvga_top (
    // Clock and reset
    .wb_clk_i	( wb_clk ),
    .wb_rst_i	( wb_rst ),
    // WISHBONE Master I/F
    .wbm_cyc_o  ( wb_vm_cyc_o ),
    .wbm_stb_o  ( wb_vm_stb_o ),
    .wbm_sel_o  ( wb_vm_sel_o ),
    .wbm_we_o   ( wb_vm_we_o ),
    .wbm_adr_o  ( wb_vm_adr_o ),
    .wbm_dat_o  ( ),
    .wbm_cab_o  ( wb_vm_cab_o ),
    .wbm_dat_i  ( wb_vm_dat_i ),
    .wbm_ack_i  ( wb_vm_ack_i ),
    .wbm_err_i  ( wb_vm_err_i ),
    .wbm_rty_i  ( 1'b0 ),
    // WISHBONE Slave I/F
    .wbs_cyc_i  ( wb_vs_cyc_i ),
    .wbs_stb_i  ( wb_vs_stb_i ),
    .wbs_sel_i  ( wb_vs_sel_i ),
    .wbs_we_i   ( wb_vs_we_i ),
    .wbs_adr_i  ( wb_vs_adr_i ),
    .wbs_dat_i  ( wb_vs_dat_i ),
    .wbs_cab_i  ( 1'b0 ),
    .wbs_dat_o  ( wb_vs_dat_o ),
    .wbs_ack_o  ( wb_vs_ack_o ),
    .wbs_err_o  ( wb_vs_err_o ),
    .wbs_rty_o  ( ),
    // Signals to VGA display
    .pad_hsync_o ( crt_hsync ),
    .pad_vsync_o ( crt_vsync ),
    .pad_rgb_o   ( {vga_r_int, vga_g_int, vga_b_int} ),
    .led_o	 ( )
);
*/
/*
CRTC_IOB crt_out_reg (
    .reset_in	( wb_rst ),
    .clk_in	( wb_clk ),
    .hsync_in	( crt_hsync ),
    .vsync_in	( crt_vsync ),
    .rgb_in	( {vga_r_int[4:1], vga_g_int[5:2], vga_b_int[4:1]} ),
    .hsync_out	( vga_hsyncn ),
    .vsync_out	( vga_vsyncn ),
    .rgb_out	( {vga_r, vga_g, vga_b} )
);
// Instantiation of the Audio controller.
// This controller connects to AK4520A Codec chip.
audio_top audio_top (
	// WISHBONE common
	.wb_clk_i ( wb_clk ),
	.wb_rst_i ( wb_rst ),
	// WISHBONE slave
	.wb_dat_i ( wb_as_dat_i ),
	.wb_adr_i ( wb_as_adr_i ),
	.wb_sel_i ( wb_as_sel_i ),
	.wb_we_i  ( wb_as_we_i  ),
	.wb_cyc_i ( wb_as_cyc_i ),
	.wb_stb_i ( wb_as_stb_i ),
	.wb_ack_o ( wb_as_ack_o ),
	.wb_err_o ( wb_as_err_o ),
	// WISHBONE master
	.m_wb_dat_o ( wb_am_dat_o ),
	.m_wb_dat_i ( wb_am_dat_i ),
	.m_wb_adr_o ( wb_am_adr_o ),
	.m_wb_sel_o ( wb_am_sel_o ),
	.m_wb_we_o  ( wb_am_we_o  ),
	.m_wb_cyc_o ( wb_am_cyc_o ),
	.m_wb_stb_o ( wb_am_stb_o ),
	.m_wb_ack_i ( wb_am_ack_i ),
	.m_wb_err_i ( wb_am_err_i ),
	// AK4520A CODEC interface
	.mclk	  ( codec_mclk ),
	.lrclk	  ( codec_lrclk ),
	.sclk	  ( codec_sclk ),
	.sdin	  ( codec_sdin ),
	.sdout	  ( codec_sdout )
);
*/
// Instantiation of the development i/f model
// Used only for simulations.
`ifdef DBG_IF_MODEL
dbg_if_model dbg_if_model  (
	// JTAG pins
	.tms_pad_i	( jtag_tms ),
	.tck_pad_i	( jtag_tck ),
	.trst_pad_i	( jtag_trst ),
	.tdi_pad_i	( jtag_tdi ),
	.tdo_pad_o	( jtag_tdo ),
	// Boundary Scan signals
	.capture_dr_o	( ),
	.shift_dr_o	( ),
	.update_dr_o	( ),
	.extest_selected_o ( ),
	.bs_chain_i	( 1'b0 ),
	// RISC signals
	.risc_clk_i	( wb_clk ),
	.risc_data_i	( dbg_dat_risc ),
	.risc_data_o	( dbg_dat_dbg ),
	.risc_addr_o	( dbg_adr ),
	.wp_i		( dbg_wp ),
	.bp_i		( dbg_bp ),
	.opselect_o	( dbg_op ),
	.lsstatus_i	( dbg_lss ),
	.istatus_i	( dbg_is ),
	.risc_stall_o	( dbg_stall ),
	.reset_o	( ),
	// WISHBONE common
	.wb_clk_i	( wb_clk ),
	.wb_rst_i	( wb_rst ),
	// WISHBONE master interface
	.wb_adr_o	( wb_dm_adr_o ),
	.wb_dat_i	( wb_dm_dat_i ),
	.wb_dat_o	( wb_dm_dat_o ),
	.wb_sel_o	( wb_dm_sel_o ),
	.wb_we_o	( wb_dm_we_o  ),
	.wb_stb_o	( wb_dm_stb_o ),
	.wb_cyc_o	( wb_dm_cyc_o ),
	.wb_cab_o	( wb_dm_cab_o ),
	.wb_ack_i	( wb_dm_ack_i ),
	.wb_err_i	( wb_dm_err_i )
);
`else
// Instantiation of the development i/f
dbg_top dbg_top  (
	// JTAG pins
	.tms_pad_i	( jtag_tms ),
	.tck_pad_i	( jtag_tck ),
	.trst_pad_i	( jtag_trst ),
	.tdi_pad_i	( jtag_tdi ),
	.tdo_pad_o	( jtag_tdo ),
	.tdo_padoen_o	( ),
	// Boundary Scan signals
	.capture_dr_o	( ),
	.shift_dr_o	( ),
	.update_dr_o	( ),
	.extest_selected_o ( ),
	.bs_chain_i	( 1'b0 ),
	.bs_chain_o	( ),
	// RISC signals
	.risc_clk_i	( wb_clk ),
	.risc_addr_o	( dbg_adr ),
	.risc_data_i	( dbg_dat_risc ),
	.risc_data_o	( dbg_dat_dbg ),
	.wp_i		( dbg_wp ),
	.bp_i		( dbg_bp ),
	.opselect_o	( dbg_op ),
	.lsstatus_i	( dbg_lss ),
	.istatus_i	( dbg_is ),
	.risc_stall_o	( dbg_stall ),
	.reset_o	( ),
	// WISHBONE common
	.wb_clk_i	( wb_clk ),
	.wb_rst_i	( wb_rst ),
	// WISHBONE master interface
	.wb_adr_o	( wb_dm_adr_o ),
	.wb_dat_i	( wb_dm_dat_i ),
	.wb_dat_o	( wb_dm_dat_o ),
	.wb_sel_o	( wb_dm_sel_o ),
	.wb_we_o	( wb_dm_we_o  ),
	.wb_stb_o	( wb_dm_stb_o ),
	.wb_cyc_o	( wb_dm_cyc_o ),
	.wb_cab_o	( wb_dm_cab_o ),
	.wb_ack_i	( wb_dm_ack_i ),
	.wb_err_i	( wb_dm_err_i )
);
`endif
// Instantiation of the OR1200 RISC
or1200_top or1200_top (
	// Common
	.rst_i		( wb_rst ),
	.clk_i		( clk ),
`ifdef OR1200_CLMODE_1TO2
	.clmode_i	( 2'b01 ),
`else
`ifdef OR1200_CLMODE_1TO4
	.clmode_i	( 2'b11 ),
`else
	.clmode_i	( 2'b00 ),
`endif
`endif
`ifdef  SPOOFER
        .clk_count      ( clk_count ),
        .spoof_out      ( spoof_out),
	.trigger	( trigger),
`endif
	// WISHBONE Instruction Master
	.iwb_clk_i	( wb_clk ),
	.iwb_rst_i	( wb_rst ),
	.iwb_cyc_o	( wb_rim_cyc_o ),
	.iwb_adr_o	( wb_rim_adr_o ),
	.iwb_dat_i	( wb_rim_dat_i ),
	.iwb_dat_o	( wb_rim_dat_o ),
	.iwb_sel_o	( wb_rim_sel_o ),
	.iwb_ack_i	( wb_rim_ack_i ),
	.iwb_err_i	( wb_rim_err_i ),
	.iwb_rty_i	( wb_rim_rty_i ),
	.iwb_we_o	( wb_rim_we_o  ),
	.iwb_stb_o	( wb_rim_stb_o ),
	.iwb_cab_o	( wb_rim_cab_o ),
	// WISHBONE Data Master
	.dwb_clk_i	( wb_clk ),
	.dwb_rst_i	( wb_rst ),
	.dwb_cyc_o	( wb_rdm_cyc_o ),
	.dwb_adr_o	( wb_rdm_adr_o ),
	.dwb_dat_i	( wb_rdm_dat_i ),
	.dwb_dat_o	( wb_rdm_dat_o ),
	.dwb_sel_o	( wb_rdm_sel_o ),
	.dwb_ack_i	( wb_rdm_ack_i ),
	.dwb_err_i	( wb_rdm_err_i ),
	.dwb_rty_i	( wb_rdm_rty_i ),
	.dwb_we_o	( wb_rdm_we_o  ),
	.dwb_stb_o	( wb_rdm_stb_o ),
	.dwb_cab_o	( wb_rdm_cab_o ),
	// Debug
	.dbg_stall_i	( dbg_stall ),
	.dbg_dat_i	( dbg_dat_dbg ),
	.dbg_adr_i	( dbg_adr ),
	.dbg_ewt_i	( 1'b0 ),
	.dbg_lss_o	( dbg_lss ),
	.dbg_is_o	( dbg_is ),
	.dbg_wp_o	( dbg_wp ),
	.dbg_bp_o	( dbg_bp ),
	.dbg_dat_o	( dbg_dat_risc ),
	.dbg_ack_o	( ),
	.dbg_stb_i	( dbg_op[2] ),
	.dbg_we_i	( dbg_op[0] ),
	// Power Management
	.pm_clksd_o	( ),
	.pm_cpustall_i	( 1'b0 ),
	.pm_dc_gate_o	( ),
	.pm_ic_gate_o	( ),
	.pm_dmmu_gate_o	( ),
	.pm_immu_gate_o	( ),
	.pm_tt_gate_o	( ),
	.pm_cpu_gate_o	( ),
	.pm_wakeup_o	( ),
	.pm_lvolt_o	( ),
	// Interrupts
	.pic_ints_i	( pic_ints )
);
// Instantiation of the Flash controller
flash_top flash_top (
	// WISHBONE common
	.wb_clk_i	( wb_clk ),
	.wb_rst_i	( wb_rst ),
	// WISHBONE slave
	.wb_dat_i	( wb_fs_dat_i ),
	.wb_dat_o	( wb_fs_dat_o ),
	.wb_adr_i	( wb_fs_adr_i ),
	.wb_sel_i	( wb_fs_sel_i ),
	.wb_we_i	( wb_fs_we_i  ),
	.wb_cyc_i	( wb_fs_cyc_i ),
	.wb_stb_i	( wb_fs_stb_i ),
	.wb_ack_o	( wb_fs_ack_o ),
	.wb_err_o	( wb_fs_err_o ),
	// Flash external
	.flash_rstn	( flash_rstn ),
	.cen		( flash_cen ),
	.oen		( flash_oen ),
	.wen		( flash_wen ),
	.rdy		( flash_rdy ),
	.d		( flash_d ),
	.a		( flash_a ),
	.a_oe		( )
);
// Instantiation of the SRAM controller
sram_top sram_top (
	// WISHBONE common
	.wb_clk_i	( wb_clk ),
	.wb_rst_i	( wb_rst ),
	// WISHBONE slave
	.wb_dat_i	( wb_ss_dat_i ),
	.wb_dat_o	( wb_ss_dat_o ),
	.wb_adr_i	( wb_ss_adr_i ),
	.wb_sel_i	( wb_ss_sel_i ),
	.wb_we_i	( wb_ss_we_i  ),
	.wb_cyc_i	( wb_ss_cyc_i ),
	.wb_stb_i	( wb_ss_stb_i ),
	.wb_ack_o	( wb_ss_ack_o ),
	.wb_err_o	( wb_ss_err_o ),
	// SRAM external
	.r_cen		( sram_r_cen ),
	.r0_wen		( sram_r0_wen ),
	.r1_wen		( sram_r1_wen ),
	.r_oen		( sram_r_oen ),
	.r_a		( sram_r_a ),
	.r_d_i		( sram_r_d ),
	.r_d_o		( sram_r_d_o ),
	.d_oe		( sram_d_oe ),
	.l_cen		( sram_l_cen ),
	.l0_wen		( sram_l0_wen ),
	.l1_wen		( sram_l1_wen ),
	.l_oen		( sram_l_oen ),
	.l_a		( sram_l_a ),
	.l_d_i		( sram_l_d ),
	.l_d_o		( sram_l_d_o )
);
// Instantiation of the UART16550
/*
uart_top uart_top (
	// WISHBONE common
	.wb_clk_i	( wb_clk ),
	.wb_rst_i	( wb_rst ),
	// WISHBONE slave
	.wb_adr_i	( wb_us_adr_i[4:0] ),
	.wb_dat_i	( wb_us_dat_i ),
	.wb_dat_o	( wb_us_dat_o ),
	.wb_we_i	( wb_us_we_i  ),
	.wb_stb_i	( wb_us_stb_i ),
	.wb_cyc_i	( wb_us_cyc_i ),
	.wb_ack_o	( wb_us_ack_o ),
	.wb_sel_i	( wb_us_sel_i ),
	// Interrupt request
	.int_o		( pic_ints[`APP_INT_UART] ),
	// UART signals
	// serial input/output
	.stx_pad_o	( uart_stx ),
	.srx_pad_i	( uart_srx ),
	// modem signals
	.rts_pad_o	( ),
	.cts_pad_i	( 1'b0 ),
	.dtr_pad_o	( ),
	.dsr_pad_i	( 1'b0 ),
	.ri_pad_i	( 1'b0 ),
	.dcd_pad_i	( 1'b0 )
);
// hdlc_ent_FCS_TYPE2_ADD_WIDTH7 hdlc_top (
hdlc_ent hdlc_top (
	// WISHBONE common
   .CLK_I    ( wb_clk ),
   .RST_I    ( wb_rst ),
	// WISHBONE slave
	.ADR_I   	( wb_hd_adr_i_map[2:0] ),
	.DAT_I	   ( wb_hd_dat_i ),
	.DAT_O	   ( wb_hd_dat_o ),
	.WE_I	    ( wb_hd_we_i ),
	.STB_I	   ( wb_hd_stb_i ),
	.CYC_I	   ( wb_hd_cyc_i ),
	.ACK_O	   ( wb_hd_ack_o ),
	.RTY_O    ( wb_hd_rty_o ),
//	.wb_sel_i	(  ),
	// Interrupt request
	.TAG0_O   ( pic_ints[`APP_INT_HDLC1] ),
	.TAG1_O   ( pic_ints[`APP_INT_HDLC2] ),
	// HDLC signals
	// serial input/output
    .Tx      ( hdlc_tx ),
    .Rx      ( hdlc_rx ),
    .Loopback ( Loopback ),
    .TxEN    ( 1'b1 ),
	 .RxEn    ( 1'b1 ),
	 .Txclk   ( tx_clk ),
	 .RxClk   ( rx_clk )
//    Txclk     : IN  STD_LOGIC;          -- Tx Clock
//    RxClk     : IN  STD_LOGIC;          -- Rx Clock
//    Tx        : OUT STD_LOGIC;          -- Tx setial line
//    Rx        : IN  STD_LOGIC;          -- Rx serial line
//    TxEN      : IN  STD_LOGIC;          -- Tx Enable
//    RxEn      : IN  STD_LOGIC;          -- Rx Enable
//    RST_I     : IN  STD_LOGIC;          -- WB reset
//    CLK_I     : IN  STD_LOGIC;          -- WB clock
//    ADR_I     : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);  -- WB address
//    DAT_O     : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);  -- WB output data
//    DAT_I     : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);  -- WB input data
//    WE_I      : IN  STD_LOGIC;          -- WB write/read signal
//    STB_I     : IN  STD_LOGIC;          -- WB strobe
//    ACK_O     : OUT STD_LOGIC;          -- WB acknowledge
//    CYC_I     : IN  STD_LOGIC;          -- WB cycle
//    RTY_O     : OUT STD_LOGIC;          -- WB Retry
//    TAG0_O    : OUT STD_LOGIC;          -- WB TAG (TxDone interrupt)
//    TAG1_O    : OUT STD_LOGIC);         -- WB TAG (RxReady interrupt)
);
*/
/*
// Instantiation of the Ethernet 10/100 MAC
eth_top eth_top (
	// WISHBONE common
	.wb_clk_i	( wb_clk ),
	.wb_rst_i	( wb_rst ),
	// WISHBONE slave
	.wb_dat_i	( wb_es_dat_i ),
	.wb_dat_o	( wb_es_dat_o ),
	.wb_adr_i	( wb_es_adr_i[11:2] ),
	.wb_sel_i	( wb_es_sel_i ),
	.wb_we_i	( wb_es_we_i  ),
	.wb_cyc_i	( wb_es_cyc_i ),
	.wb_stb_i	( wb_es_stb_i ),
	.wb_ack_o	( wb_es_ack_o ),
	.wb_err_o	( wb_es_err_o ),
	// WISHBONE master
	.m_wb_adr_o	( wb_em_adr_o ),
	.m_wb_sel_o	( wb_em_sel_o ),
	.m_wb_we_o	( wb_em_we_o  ),
	.m_wb_dat_o	( wb_em_dat_o ),
	.m_wb_dat_i	( wb_em_dat_i ),
	.m_wb_cyc_o	( wb_em_cyc_o ),
	.m_wb_stb_o	( wb_em_stb_o ),
	.m_wb_ack_i	( wb_em_ack_i ),
	.m_wb_err_i	( wb_em_err_i ),
	// TX
	.mtx_clk_pad_i	( eth_tx_clk ),
	.mtxd_pad_o	( eth_txd ),
	.mtxen_pad_o	( eth_tx_en ),
	.mtxerr_pad_o	( eth_tx_er ),
	// RX
	.mrx_clk_pad_i	( eth_rx_clk ),
	.mrxd_pad_i	( eth_rxd ),
	.mrxdv_pad_i	( eth_rx_dv ),
	.mrxerr_pad_i	( eth_rx_er ),
	.mcoll_pad_i	( eth_col ),
	.mcrs_pad_i	( eth_crs ),
	// MIIM
	.mdc_pad_o	( eth_mdc ),
	.md_pad_i	( eth_mdio ),
	.md_pad_o	( eth_mdo ),
	.md_padoe_o	( eth_mdoe ),
	// Interrupt
	.int_o		( pic_ints[`APP_INT_ETH] )
);
*/
/*
// Instantiation of the PS/2 Keyboard Controller
ps2_top ps2_top (
	// WISHBONE common
	.wb_clk_i	( wb_clk ),
	.wb_rst_i	( wb_rst ),
	// WISHBONE slave
	.wb_cyc_i	( wb_ps_cyc_i ),
	.wb_stb_i	( wb_ps_stb_i ),
	.wb_we_i	( wb_ps_we_i  ),
	.wb_sel_i	( wb_ps_sel_i ),
	.wb_adr_i	( wb_ps_adr_i ),
	.wb_dat_i	( wb_ps_dat_i ),
	.wb_dat_o	( wb_ps_dat_o ),
	.wb_ack_o	( wb_ps_ack_o ),
	// Interrupt
	.wb_int_o	( pic_ints[`APP_INT_PS2] ),
	// PS/2 external wires
	.ps2_kbd_clk_pad_i	( ps2_clk ),
	.ps2_kbd_data_pad_i	( ps2_data ),
	.ps2_kbd_clk_pad_o	( ps2_clk_o ),
	.ps2_kbd_data_pad_o	( ps2_data_o ),
	.ps2_kbd_clk_pad_oe_o	( ps2_clk_oe ),
	.ps2_kbd_data_pad_oe_o	( ps2_data_oe )
);
*/
// Instantiation of the CPLD TDM
// This small block connects XSV FPGA (xsv_fpga_top)
// to the CPLD. CPLD has connections to the
// RS232 PHY chip and to host PC (if you run OR1K
// GDB debugger). In order for TDM to work, CPLD
// must also be programmed with TDM master i/f.
tdm_slave_if tdm_slave_if (
	.clk	( wb_clk ),
	.rst	( wb_rst ),
	.tdmfrm	( tdmfrm ),
	.tdmrx	( tdmrx ),
	.tdmtx	( tdmtx ),
	.din	( { jtag_tdo, uart_stx, 6'b000_000 } ),
	.dout	( { jtag_tms, jtag_tck, jtag_trst, jtag_tdi, uart_srx, tdm_out_unused } )
);
// Instantiation of the Traffic COP
tc_top #(`APP_ADDR_DEC_W,
	 `APP_ADDR_SRAM,
	 `APP_ADDR_DEC_W,
	 `APP_ADDR_FLASH,
	 `APP_ADDR_DECP_W,
	 `APP_ADDR_PERIP,
	 `APP_ADDR_DEC_W,
	 `APP_ADDR_VGA,
	 `APP_ADDR_ETH,
	 `APP_ADDR_AUDIO,
//	 `APP_ADDR_UART,
//	 `APP_ADDR_PS2,
//	 `APP_ADDR_HDLC,
	 `APP_ADDR_RES2
	) tc_top (
	// WISHBONE common
	.wb_clk_i	( wb_clk ),
	.wb_rst_i	( wb_rst ),
	// WISHBONE Initiator 0
	/*
	.i0_wb_cyc_i	( wb_vm_cyc_o ),
	.i0_wb_stb_i	( wb_vm_stb_o ),
	.i0_wb_cab_i	( wb_vm_cab_o ),
	.i0_wb_adr_i	( wb_vm_adr_o ),
	.i0_wb_sel_i	( wb_vm_sel_o ),
	.i0_wb_we_i	( wb_vm_we_o  ),
	.i0_wb_dat_i	( 32'h0000_0000 ),
	.i0_wb_dat_o	( wb_vm_dat_i ),
	.i0_wb_ack_o	( wb_vm_ack_i ),
	.i0_wb_err_o	( wb_vm_err_i ),
	.i0_wb_cyc_i	( 1'b0 ),
	.i0_wb_stb_i	( 1'b0 ),
	.i0_wb_cab_i	( 1'b0 ),
	.i0_wb_adr_i	( 32'h0000_0000 ),
	.i0_wb_sel_i	( 4'b0000 ),
	.i0_wb_we_i	( 1'b0 ),
	.i0_wb_dat_i	( 32'h0000_0000 ),
	.i0_wb_dat_o	( ),
	.i0_wb_ack_o	( ),
	.i0_wb_err_o	( ),
	// WISHBONE Initiator 1
	.i0_wb_cyc_i	( wb_em_cyc_o ),
	.i0_wb_stb_i	( wb_em_stb_o ),
	.i0_wb_cab_i	( wb_em_cab_o ),
	.i0_wb_adr_i	( wb_em_adr_o ),
	.i0_wb_sel_i	( wb_em_sel_o ),
	.i0_wb_we_i	( wb_em_we_o  ),
	.i0_wb_dat_i	( wb_em_dat_o ),
	.i0_wb_dat_o	( wb_em_dat_i ),
	.i0_wb_ack_o	( wb_em_ack_i ),
	.i0_wb_err_o	( wb_em_err_i ),
	// WISHBONE Initiator 2
	.i1_wb_cyc_i	( wb_am_cyc_o ),
	.i1_wb_stb_i	( wb_am_stb_o ),
	.i1_wb_cab_i	( wb_am_cab_o ),
	.i1_wb_adr_i	( wb_am_adr_o ),
	.i1_wb_sel_i	( wb_am_sel_o ),
	.i1_wb_we_i	( wb_am_we_o  ),
	.i1_wb_dat_i	( wb_am_dat_o ),
	.i1_wb_dat_o	( wb_am_dat_i ),
	.i1_wb_ack_o	( wb_am_ack_i ),
	.i1_wb_err_o	( wb_am_err_i ),
	// WISHBONE Initiator 3
	.i3_wb_cyc_i	( wb_dm_cyc_o ),
	.i3_wb_stb_i	( wb_dm_stb_o ),
	.i3_wb_cab_i	( wb_dm_cab_o ),
	.i3_wb_adr_i	( wb_dm_adr_o ),
	.i3_wb_sel_i	( wb_dm_sel_o ),
	.i3_wb_we_i	( wb_dm_we_o  ),
	.i3_wb_dat_i	( wb_dm_dat_o ),
	.i3_wb_dat_o	( wb_dm_dat_i ),
	.i3_wb_ack_o	( wb_dm_ack_i ),
	.i3_wb_err_o	( wb_dm_err_i ),
*/
	.i0_wb_cyc_i	( 1'b0 ),
	.i0_wb_stb_i	( 1'b0 ),
	.i0_wb_cab_i	( 1'b0 ),
	.i0_wb_adr_i	( 32'h0000_0000 ),
	.i0_wb_sel_i	( 4'b0000 ),
	.i0_wb_we_i	( 1'b0 ),
	.i0_wb_dat_i	( 32'h0000_0000 ),
	.i0_wb_dat_o	( ),
	.i0_wb_ack_o	( ),
	.i0_wb_err_o	( ),
	.i1_wb_cyc_i	( 1'b0 ),
	.i1_wb_stb_i	( 1'b0 ),
	.i1_wb_cab_i	( 1'b0 ),
	.i1_wb_adr_i	( 32'h0000_0000 ),
	.i1_wb_sel_i	( 4'b0000 ),
	.i1_wb_we_i	( 1'b0 ),
	.i1_wb_dat_i	( 32'h0000_0000 ),
	.i1_wb_dat_o	( ),
	.i1_wb_ack_o	( ),
	.i1_wb_err_o	( ),
	.i2_wb_cyc_i	( 1'b0 ),
	.i2_wb_stb_i	( 1'b0 ),
	.i2_wb_cab_i	( 1'b0 ),
	.i2_wb_adr_i	( 32'h0000_0000 ),
	.i2_wb_sel_i	( 4'b0000 ),
	.i2_wb_we_i	( 1'b0 ),
	.i2_wb_dat_i	( 32'h0000_0000 ),
	.i2_wb_dat_o	( ),
	.i2_wb_ack_o	( ),
	.i2_wb_err_o	( ),
	.i3_wb_cyc_i	( 1'b0 ),
	.i3_wb_stb_i	( 1'b0 ),
	.i3_wb_cab_i	( 1'b0 ),
	.i3_wb_adr_i	( 32'h0000_0000 ),
	.i3_wb_sel_i	( 4'b0000 ),
	.i3_wb_we_i	( 1'b0 ),
	.i3_wb_dat_i	( 32'h0000_0000 ),
	.i3_wb_dat_o	( ),
	.i3_wb_ack_o	( ),
	.i3_wb_err_o	( ),
	// WISHBONE Initiator 4
	.i4_wb_cyc_i	( wb_rdm_cyc_o ),
	.i4_wb_stb_i	( wb_rdm_stb_o ),
	.i4_wb_cab_i	( wb_rdm_cab_o ),
	.i4_wb_adr_i	( wb_rdm_adr_o ),
	.i4_wb_sel_i	( wb_rdm_sel_o ),
	.i4_wb_we_i	( wb_rdm_we_o  ),
	.i4_wb_dat_i	( wb_rdm_dat_o ),
	.i4_wb_dat_o	( wb_rdm_dat_i ),
	.i4_wb_ack_o	( wb_rdm_ack ),
	.i4_wb_err_o	( wb_rdm_err_i ),
	// WISHBONE Initiator 5
	.i5_wb_cyc_i	( wb_rim_cyc_o ),
	.i5_wb_stb_i	( wb_rim_stb_o ),
	.i5_wb_cab_i	( wb_rim_cab_o ),
	.i5_wb_adr_i	( wb_rif_adr ),
	.i5_wb_sel_i	( wb_rim_sel_o ),
	.i5_wb_we_i	( wb_rim_we_o  ),
	.i5_wb_dat_i	( wb_rim_dat_o ),
	.i5_wb_dat_o	( wb_rim_dat_i ),
	.i5_wb_ack_o	( wb_rim_ack_i ),
	.i5_wb_err_o	( wb_rim_err_i ),
	// WISHBONE Initiator 6
	.i6_wb_cyc_i	( 1'b0 ),
	.i6_wb_stb_i	( 1'b0 ),
	.i6_wb_cab_i	( 1'b0 ),
	.i6_wb_adr_i	( 32'h0000_0000 ),
	.i6_wb_sel_i	( 4'b0000 ),
	.i6_wb_we_i	( 1'b0 ),
	.i6_wb_dat_i	( 32'h0000_0000 ),
	.i6_wb_dat_o	( ),
	.i6_wb_ack_o	( ),
	.i6_wb_err_o	( ),
	// WISHBONE Initiator 7
	.i7_wb_cyc_i	( 1'b0 ),
	.i7_wb_stb_i	( 1'b0 ),
	.i7_wb_cab_i	( 1'b0 ),
	.i7_wb_adr_i	( 32'h0000_0000 ),
	.i7_wb_sel_i	( 4'b0000 ),
	.i7_wb_we_i	( 1'b0 ),
	.i7_wb_dat_i	( 32'h0000_0000 ),
	.i7_wb_dat_o	( ),
	.i7_wb_ack_o	( ),
	.i7_wb_err_o	( ),
	// WISHBONE Target 0
	.t0_wb_cyc_o	( wb_ss_cyc_i ),
	.t0_wb_stb_o	( wb_ss_stb_i ),
	.t0_wb_cab_o	( wb_ss_cab_i ),
	.t0_wb_adr_o	( wb_ss_adr_i ),
	.t0_wb_sel_o	( wb_ss_sel_i ),
	.t0_wb_we_o	( wb_ss_we_i  ),
	.t0_wb_dat_o	( wb_ss_dat_i ),
	.t0_wb_dat_i	( wb_ss_dat_o ),
	.t0_wb_ack_i	( wb_ss_ack_o ),
	.t0_wb_err_i	( wb_ss_err_o ),
	// WISHBONE Target 1
	.t1_wb_cyc_o	( wb_fs_cyc_i ),
	.t1_wb_stb_o	( wb_fs_stb_i ),
	.t1_wb_cab_o	( wb_fs_cab_i ),
	.t1_wb_adr_o	( wb_fs_adr_i ),
	.t1_wb_sel_o	( wb_fs_sel_i ),
	.t1_wb_we_o	( wb_fs_we_i  ),
	.t1_wb_dat_o	( wb_fs_dat_i ),
	.t1_wb_dat_i	( wb_fs_dat_o ),
	.t1_wb_ack_i	( wb_fs_ack_o ),
	.t1_wb_err_i	( wb_fs_err_o ),
	.t2_wb_cyc_o	( ),
	.t2_wb_stb_o	( ),
	.t2_wb_cab_o	( ),
	.t2_wb_adr_o	( ),
	.t2_wb_sel_o	( ),
	.t2_wb_we_o	( ),
	.t2_wb_dat_o	( ),
	.t2_wb_dat_i	( 32'h0000_0000 ),
	.t2_wb_ack_i	( 1'b0 ),
	.t2_wb_err_i	( 1'b1 ),
	.t3_wb_cyc_o	( ),
	.t3_wb_stb_o	( ),
	.t3_wb_cab_o	( ),
	.t3_wb_adr_o	( ),
	.t3_wb_sel_o	( ),
	.t3_wb_we_o	( ),
	.t3_wb_dat_o	( ),
	.t3_wb_dat_i	( 32'h0000_0000 ),
	.t3_wb_ack_i	( 1'b0 ),
	.t3_wb_err_i	( 1'b1 ),
	.t4_wb_cyc_o	( ),
	.t4_wb_stb_o	( ),
	.t4_wb_cab_o	( ),
	.t4_wb_adr_o	( ),
	.t4_wb_sel_o	( ),
	.t4_wb_we_o	( ),
	.t4_wb_dat_o	( ),
	.t4_wb_dat_i	( 32'h0000_0000 ),
	.t4_wb_ack_i	( 1'b0 ),
	.t4_wb_err_i	( 1'b1 ),
	.t5_wb_cyc_o	( ),
	.t5_wb_stb_o	( ),
	.t5_wb_cab_o	( ),
	.t5_wb_adr_o	( ),
	.t5_wb_sel_o	( ),
	.t5_wb_we_o	( ),
	.t5_wb_dat_o	( ),
	.t5_wb_dat_i	( 32'h0000_0000 ),
	.t5_wb_ack_i	( 1'b0 ),
	.t5_wb_err_i	( 1'b1 ),
	.t6_wb_cyc_o	( ),
	.t6_wb_stb_o	( ),
	.t6_wb_cab_o	( ),
	.t6_wb_adr_o	( ),
	.t6_wb_sel_o	( ),
	.t6_wb_we_o	( ),
	.t6_wb_dat_o	( ),
	.t6_wb_dat_i	( 32'h0000_0000 ),
	.t6_wb_ack_i	( 1'b0 ),
	.t6_wb_err_i	( 1'b1 ),
	.t7_wb_cyc_o	( ),
	.t7_wb_stb_o	( ),
	.t7_wb_cab_o	( ),
	.t7_wb_adr_o	( ),
	.t7_wb_sel_o	( ),
	.t7_wb_we_o	( ),
	.t7_wb_dat_o	( ),
	.t7_wb_dat_i	( 32'h0000_0000 ),
	.t7_wb_ack_i	( 1'b0 ),
	.t7_wb_err_i	( 1'b1 ),
        /*
        // WISHBONE Target 2
	.t2_wb_cyc_o	( wb_vs_cyc_i ),
	.t2_wb_stb_o	( wb_vs_stb_i ),
	.t2_wb_cab_o	( wb_vs_cab_i ),
	.t2_wb_adr_o	( wb_vs_adr_i ),
	.t2_wb_sel_o	( wb_vs_sel_i ),
	.t2_wb_we_o	( wb_vs_we_i  ),
	.t2_wb_dat_o	( wb_vs_dat_i ),
	.t2_wb_dat_i	( wb_vs_dat_o ),
	.t2_wb_ack_i	( wb_vs_ack_o ),
	.t2_wb_err_i	( wb_vs_err_o ),
	// WISHBONE Target 3
	.t3_wb_cyc_o	( wb_es_cyc_i ),
	.t3_wb_stb_o	( wb_es_stb_i ),
	.t3_wb_cab_o	( wb_es_cab_i ),
	.t3_wb_adr_o	( wb_es_adr_i ),
	.t3_wb_sel_o	( wb_es_sel_i ),
	.t3_wb_we_o	( wb_es_we_i  ),
	.t3_wb_dat_o	( wb_es_dat_i ),
	.t3_wb_dat_i	( wb_es_dat_o ),
	.t3_wb_ack_i	( wb_es_ack_o ),
	.t3_wb_err_i	( wb_es_err_o ),
	// WISHBONE Target 4
	.t4_wb_cyc_o	( wb_as_cyc_i ),
	.t4_wb_stb_o	( wb_as_stb_i ),
	.t4_wb_cab_o	( wb_as_cab_i ),
	.t4_wb_adr_o	( wb_as_adr_i ),
	.t4_wb_sel_o	( wb_as_sel_i ),
	.t4_wb_we_o	( wb_as_we_i  ),
	.t4_wb_dat_o	( wb_as_dat_i ),
	.t4_wb_dat_i	( wb_as_dat_o ),
	.t4_wb_ack_i	( wb_as_ack_o ),
	.t4_wb_err_i	( wb_as_err_o ),
	// WISHBONE Target 5
	.t5_wb_cyc_o	( wb_us_cyc_i ),
	.t5_wb_stb_o	( wb_us_stb_i ),
	.t5_wb_cab_o	( wb_us_cab_i ),
	.t5_wb_adr_o	( wb_us_adr_i ),
	.t5_wb_sel_o	( wb_us_sel_i ),
	.t5_wb_we_o	( wb_us_we_i  ),
	.t5_wb_dat_o	( wb_us_dat_i ),
	.t5_wb_dat_i	( wb_us_dat_o ),
	.t5_wb_ack_i	( wb_us_ack_o ),
	.t5_wb_err_i	( wb_us_err_o ),
	// WISHBONE Target 6
	.t6_wb_cyc_o	( wb_ps_cyc_i ),
	.t6_wb_stb_o	( wb_ps_stb_i ),
	.t6_wb_cab_o	( wb_ps_cab_i ),
	.t6_wb_adr_o	( wb_ps_adr_i ),
	.t6_wb_sel_o	( wb_ps_sel_i ),
	.t6_wb_we_o	( wb_ps_we_i  ),
	.t6_wb_dat_o	( wb_ps_dat_i ),
	.t6_wb_dat_i	( wb_ps_dat_o ),
	.t6_wb_ack_i	( wb_ps_ack_o ),
	.t6_wb_err_i	( wb_ps_err_o ),
	// WISHBONE Target 7
	.t7_wb_cyc_o	( wb_hd_cyc_i ),
	.t7_wb_stb_o	( wb_hd_stb_i ),
	.t7_wb_cab_o	( wb_hd_cab_i ),
	.t7_wb_adr_o	( wb_hd_adr_i ),
	.t7_wb_sel_o	( wb_hd_sel_i ),
	.t7_wb_we_o	 ( wb_hd_we_i  ),
	.t7_wb_dat_o	( wb_hd_dat_i ),
	.t7_wb_dat_i	( wb_hd_dat_o ),
	.t7_wb_ack_i	( wb_hd_ack_o ),
	.t7_wb_err_i	( wb_hd_err_o ),
        */
	// WISHBONE Target 8
	.t8_wb_cyc_o	( ),
	.t8_wb_stb_o	( ),
	.t8_wb_cab_o	( ),
	.t8_wb_adr_o	( ),
	.t8_wb_sel_o	( ),
	.t8_wb_we_o	( ),
	.t8_wb_dat_o	( ),
	.t8_wb_dat_i	( 32'h0000_0000 ),
	.t8_wb_ack_i	( 1'b0 ),
	.t8_wb_err_i	( 1'b1 )
);
//initial begin
//  $dumpvars(0);
//  $dumpfile("dump.vcd");
//end
endmodule