module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_a
		inst_a_e inst_a (
		);
		// End of Generated Instance Port Map for inst_a
		// Generated Instance Port Map for inst_e
		inst_e_e inst_e (
		);
		// End of Generated Instance Port Map for inst_e
endmodule