module  rg66dae (
   sys_clk,
   rst_n,
   ls35987,
   yzae707,
   fa7383c,
   ng9c1e2,
   qge0f13,
   qv7898,
   an3c4c4,
   ene2624,
   zz13124,
   aa98926,
   mec4930,
   wy24981,
   ks24c08,
   wwf5804,
   vk30204,
   wyac021,
   uv60109,
   ym84d,
   pu4269,
   qi2134a,
   bn169d7,
   wlb4ebf,
   xya75fd
   );
parameter  tw3afea = 1'b0;
parameter  bld7f52  = 1'b1;
input                     sys_clk;
input                     rst_n;
input                     ls35987;
input  [15:0]             yzae707;
input                     fa7383c;
input                     ng9c1e2;
input                     qge0f13;
input                     qv7898;
input                     an3c4c4;
input                     ene2624;
input                     zz13124;
input                     aa98926;
input                     wy24981;
input  [15:0]             ks24c08;
input  [3:0]              mec4930;
output [15:0]             wwf5804;
output                    vk30204;
output                    wyac021;
output                    uv60109;
output                    ym84d;
output                    pu4269;
output                    qi2134a;
output                    bn169d7;
output                    wlb4ebf;
output                    xya75fd;
reg    [15:0]             wwf5804;
reg                       vk30204;
reg                       wyac021;
reg                       uv60109;
reg                       ym84d;
reg                       pu4269;
reg                       qi2134a;
reg                       bn169d7;
reg                       wlb4ebf;
reg                       xya75fd;
reg    [15:0]             mt295f, tw14afc, hda57e2, czf8578, vvc2bc4, mg15e26, dbaf130, su78986;
reg                       uic4c31;
reg                       kf26189,  tw30c4c,  zm86263,  wy3131b,  tw898d8,  ea4c6c3,  lq63618, ba1b0c2;
reg                       xjd8612,    uvc3097,    kf184bd,    vvc25ed,    sj12f6f,    aa97b7d,    ngbdbe9,   ipedf4b;
reg                       ip6fa5c,   kq7d2e5,   hbe9728,   en4b947,   kq5ca3c,   ose51e0,   fp28f01,  jc4780e;
reg                       wl3c072,   wwe0394,   pu1ca1,   vke50b,   ui7285b,   fp942d8,   cba16c7,  lsb63d;
reg                       uv5b1eb, thd8f5c, ldc7ae6, nt3d736;
reg                       dmeb9b6;
reg  [3:0]                ww5cdb3;
reg  [1:0]                jpe6d98;
reg  [7:0]                qv36cc7;
reg bl64b01;
reg [15 : 0] wyb31e1;
reg wy98f09;
reg jpc7848;
reg wl3c246;
reg xwe1234;
reg zz91a3;
reg xw48d1e;
reg kq468f3;
reg co34798;
reg [3 : 0] oua3cc0;
reg do1e601;
reg [15 : 0] nrf300a;
reg [15 : 0] ld64bcd;
reg [15 : 0] ba25e6e;
reg [15 : 0] zm2f372;
reg [15 : 0] ouae52;
reg [15 : 0] ne57290;
reg [15 : 0] ieb9482;
reg [15 : 0] psca410;
reg [15 : 0] zk52083;
reg cb9041a;
reg co820d5;
reg uk106a9;
reg ri83549;
reg ks1aa4b;
reg tud5259;
reg iea92cb;
reg kq49659;
reg ip4b2c8;
reg ui59645;
reg uicb229;
reg me59149;
reg ldc8a49;
reg vv4524f;
reg oh2927e;
reg go493f5;
reg ay49fa8;
reg ld4fd41;
reg rt7ea0e;
reg icf5076;
reg lsa83b0;
reg kd41d83;
reg hqec1d;
reg jc760ea;
reg zzb0753;
reg ri83a9e;
reg ir1d4f2;
reg cmea795;
reg kq53ca8;
reg rv9e541;
reg uvf2a0e;
reg ep95074;
reg twa83a5;
reg wj41d2b;
reg zme95d;
reg zx74aea;
reg xla5757;
reg wy2babf;
reg [3 : 0] tu5d5f9;
reg [1 : 0] meeafcb;
reg [7 : 0] rg57e59;
reg [2047:0] necf6c2;
wire [61:0] ld7b613;
localparam qgdb09f = 62,nrd84f8 = 32'hfdffd84b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      uic4c31  <= 1'b0;      mt295f <= 0; kf26189  <= 1'b0; xjd8612    <= 1'b0; ip6fa5c   <= 1'b0; wl3c072   <= 1'b0;      tw14afc <= 0; tw30c4c  <= 1'b0; uvc3097    <= 1'b0; kq7d2e5   <= 1'b0; wwe0394   <= 1'b0;      hda57e2 <= 0; zm86263  <= 1'b0; kf184bd    <= 1'b0; hbe9728   <= 1'b0; pu1ca1   <= 1'b0;      czf8578 <= 0; wy3131b  <= 1'b0; vvc25ed    <= 1'b0; en4b947   <= 1'b0; vke50b   <= 1'b0;      vvc2bc4 <= 0; tw898d8  <= 1'b0; sj12f6f    <= 1'b0; kq5ca3c   <= 1'b0; ui7285b   <= 1'b0;      mg15e26 <= 0; ea4c6c3  <= 1'b0; aa97b7d    <= 1'b0; ose51e0   <= 1'b0; fp942d8   <= 1'b0;      dbaf130 <= 0; lq63618  <= 1'b0; ngbdbe9    <= 1'b0; fp28f01   <= 1'b0; cba16c7   <= 1'b0;      su78986 <= 0; ba1b0c2  <= 1'b0; ipedf4b    <= 1'b0; jc4780e   <= 1'b0; lsb63d   <= 1'b0;   end   else begin      uic4c31  <= wy98f09;      mt295f <= wyb31e1; kf26189 <= cb9041a; xjd8612 <= jpc7848; ip6fa5c <= wl3c246; wl3c072 <= xwe1234;      tw14afc <= ld64bcd;     tw30c4c <= co820d5;     uvc3097 <= ui59645;     kq7d2e5 <= ld4fd41;     wwe0394 <= ri83a9e;      hda57e2 <= ba25e6e;     zm86263 <= uk106a9;     kf184bd <= uicb229;     hbe9728 <= rt7ea0e;     pu1ca1 <= ir1d4f2;      czf8578 <= zm2f372;     wy3131b <= ri83549;     vvc25ed <= me59149;     en4b947 <= icf5076;     vke50b <= cmea795;      vvc2bc4 <= ouae52;     tw898d8 <= ks1aa4b;     sj12f6f <= ldc8a49;     kq5ca3c <= lsa83b0;     ui7285b <= kq53ca8;      mg15e26 <= ne57290;     ea4c6c3 <= tud5259;     aa97b7d <= vv4524f;     ose51e0 <= kd41d83;     fp942d8 <= rv9e541;      dbaf130 <= ieb9482;     lq63618 <= iea92cb;     ngbdbe9 <= oh2927e;     fp28f01 <= hqec1d;     cba16c7 <= uvf2a0e;      su78986 <= psca410;     ba1b0c2 <= kq49659;     ipedf4b <= go493f5;     jc4780e <= jc760ea;     lsb63d <= ep95074;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      wwf5804     <= 0;      vk30204      <= 1'b0;      wyac021       <= 1'b0;      uv60109      <= 1'b0;      ym84d      <= 1'b0;      pu4269  <= 1'b0;      qi2134a <= 1'b0;      bn169d7     <= 1'b0;      qv36cc7    <= 8'h00;   end   else begin      pu4269     <= kq468f3;      qi2134a    <= co34798;      qv36cc7       <= nrf300a[7:0];            bn169d7        <= xla5757;            wwf5804        <= do1e601 ? {rg57e59, nrf300a[15:8]} : {zk52083[7:0], psca410[15:8]};      vk30204         <= kq49659 | do1e601 | xla5757;      wyac021          <= go493f5;                  uv60109         <= zzb0753;      ym84d         <= twa83a5;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      dmeb9b6    <= tw3afea;      wlb4ebf     <= 1'b0;      xya75fd     <= 1'b0;      jpe6d98       <= 2'b00;      ww5cdb3 <= 4'b0000;      uv5b1eb     <= 1'b0;      thd8f5c    <= 1'b0;      ldc7ae6    <= 1'b0;      nt3d736    <= 1'b0;   end   else begin      thd8f5c  <= wj41d2b;      ldc7ae6  <= zme95d;      nt3d736  <= zx74aea;                        case(wy2babf)         tw3afea : begin                         uv5b1eb  <= 1'b0;            wlb4ebf  <= 1'b0;            xya75fd  <= 1'b0;            jpe6d98    <= 2'b00;            if(!cb9041a && !co820d5 && !uk106a9 && !ri83549 && !ks1aa4b) begin                if(oua3cc0 != tu5d5f9) begin                  dmeb9b6    <= bld7f52;                  uv5b1eb     <= 1'b1;                  ww5cdb3 <= tu5d5f9 + 4'd1;               end               else if(zz91a3) begin                  dmeb9b6    <= bld7f52;                  wlb4ebf     <= 1'b1;                  xya75fd     <= 1'b0;               end               else if(xw48d1e) begin                  dmeb9b6    <= bld7f52;                  wlb4ebf     <= 1'b0;                  xya75fd     <= 1'b1;               end            end         end         bld7f52 : begin            wlb4ebf  <= 1'b0;            xya75fd  <= 1'b0;            jpe6d98    <= meeafcb + 1'b1;                                    if(wj41d2b)               dmeb9b6  <= tw3afea;            else if(meeafcb == 2'b10)               dmeb9b6  <= tw3afea;         end         default : begin            dmeb9b6    <= tw3afea;         end      endcase   end
end
always@* begin bl64b01<=ld7b613[0];wyb31e1<={yzae707>>1,ld7b613[1]};wy98f09<=ld7b613[2];jpc7848<=ld7b613[3];wl3c246<=ld7b613[4];xwe1234<=ld7b613[5];zz91a3<=ld7b613[6];xw48d1e<=ld7b613[7];kq468f3<=ld7b613[8];co34798<=ld7b613[9];oua3cc0<={mec4930>>1,ld7b613[10]};do1e601<=ld7b613[11];nrf300a<={ks24c08>>1,ld7b613[12]};ld64bcd<={mt295f>>1,ld7b613[13]};ba25e6e<={tw14afc>>1,ld7b613[14]};zm2f372<={hda57e2>>1,ld7b613[15]};ouae52<={czf8578>>1,ld7b613[16]};ne57290<={vvc2bc4>>1,ld7b613[17]};ieb9482<={mg15e26>>1,ld7b613[18]};psca410<={dbaf130>>1,ld7b613[19]};zk52083<={su78986>>1,ld7b613[20]};cb9041a<=ld7b613[21];co820d5<=ld7b613[22];uk106a9<=ld7b613[23];ri83549<=ld7b613[24];ks1aa4b<=ld7b613[25];tud5259<=ld7b613[26];iea92cb<=ld7b613[27];kq49659<=ld7b613[28];ip4b2c8<=ld7b613[29];ui59645<=ld7b613[30];uicb229<=ld7b613[31];me59149<=ld7b613[32];ldc8a49<=ld7b613[33];vv4524f<=ld7b613[34];oh2927e<=ld7b613[35];go493f5<=ld7b613[36];ay49fa8<=ld7b613[37];ld4fd41<=ld7b613[38];rt7ea0e<=ld7b613[39];icf5076<=ld7b613[40];lsa83b0<=ld7b613[41];kd41d83<=ld7b613[42];hqec1d<=ld7b613[43];jc760ea<=ld7b613[44];zzb0753<=ld7b613[45];ri83a9e<=ld7b613[46];ir1d4f2<=ld7b613[47];cmea795<=ld7b613[48];kq53ca8<=ld7b613[49];rv9e541<=ld7b613[50];uvf2a0e<=ld7b613[51];ep95074<=ld7b613[52];twa83a5<=ld7b613[53];wj41d2b<=ld7b613[54];zme95d<=ld7b613[55];zx74aea<=ld7b613[56];xla5757<=ld7b613[57];wy2babf<=ld7b613[58];tu5d5f9<={ww5cdb3>>1,ld7b613[59]};meeafcb<={jpe6d98>>1,ld7b613[60]};rg57e59<={qv36cc7>>1,ld7b613[61]};end
always@* begin necf6c2[2047]<=yzae707[0];necf6c2[2046]<=fa7383c;necf6c2[2044]<=ng9c1e2;necf6c2[2040]<=qge0f13;necf6c2[2033]<=qv7898;necf6c2[2019]<=an3c4c4;necf6c2[1999]<=aa97b7d;necf6c2[1991]<=ene2624;necf6c2[1981]<=fp942d8;necf6c2[1958]<=ldc7ae6;necf6c2[1950]<=ngbdbe9;necf6c2[1947]<=kq5ca3c;necf6c2[1934]<=zz13124;necf6c2[1914]<=cba16c7;necf6c2[1892]<=su78986[0];necf6c2[1868]<=nt3d736;necf6c2[1852]<=ipedf4b;necf6c2[1851]<=hda57e2[0];necf6c2[1847]<=ose51e0;necf6c2[1820]<=aa98926;necf6c2[1783]<=pu1ca1;necf6c2[1780]<=lsb63d;necf6c2[1737]<=uic4c31;necf6c2[1689]<=dmeb9b6;necf6c2[1657]<=ip6fa5c;necf6c2[1654]<=czf8578[0];necf6c2[1647]<=fp28f01;necf6c2[1610]<=zm86263;necf6c2[1593]<=mec4930[0];necf6c2[1523]<=vvc25ed;necf6c2[1519]<=vke50b;necf6c2[1513]<=uv5b1eb;necf6c2[1426]<=kf26189;necf6c2[1404]<=uvc3097;necf6c2[1330]<=ww5cdb3[0];necf6c2[1267]<=kq7d2e5;necf6c2[1260]<=vvc2bc4[0];necf6c2[1246]<=jc4780e;necf6c2[1225]<=qv36cc7[0];necf6c2[1199]<=lq63618;necf6c2[1173]<=wy3131b;necf6c2[1139]<=wy24981;necf6c2[1023]<=ls35987;necf6c2[999]<=sj12f6f;necf6c2[990]<=ui7285b;necf6c2[979]<=thd8f5c;necf6c2[973]<=en4b947;necf6c2[946]<=dbaf130[0];necf6c2[925]<=tw14afc[0];necf6c2[891]<=wwe0394;necf6c2[805]<=tw30c4c;necf6c2[761]<=kf184bd;necf6c2[702]<=xjd8612;necf6c2[612]<=jpe6d98[0];necf6c2[599]<=ea4c6c3;necf6c2[486]<=hbe9728;necf6c2[473]<=mg15e26[0];necf6c2[462]<=mt295f[0];necf6c2[445]<=wl3c072;necf6c2[351]<=ba1b0c2;necf6c2[299]<=tw898d8;necf6c2[231]<=ks24c08[0];end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule