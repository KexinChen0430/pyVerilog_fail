module to test
    min_max_tracker tracker(clk, adc_d, 8'd127, min, max);
endmodule