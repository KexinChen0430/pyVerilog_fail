module matchfilter_st (clk,
              rst,
              data_in,
              clk_en,
              rdy_to_ld,
              done,
              fir_result);
parameter DATA_WIDTH  = 15;
parameter COEF_WIDTH  = 13;
parameter ACCUM_WIDTH = 31;
parameter MSB_RM = 0;
parameter LSB_RM = 1;
parameter WIDTH_SAT = ACCUM_WIDTH-LSB_RM;
input clk, rst;
input [DATA_WIDTH-1:0] data_in;
input clk_en;
output rdy_to_ld;
wire rdy_to_ld;
wire rdy_int;
wire data_ld;
output done;
wire done;
wire done_int;
output [ACCUM_WIDTH-MSB_RM-LSB_RM-1:0] fir_result;
wire addr_low;
assign addr_low = 1'b0;
wire inv_rst;
assign inv_rst = ~rst;
assign data_ld = rdy_int;
wire [14:0] tdl_0_n;
wire [14:0] tdl_1_n;
wire [14:0] tdl_2_n;
wire [14:0] tdl_3_n;
wire [14:0] tdl_4_n;
wire [14:0] tdl_5_n;
wire [14:0] tdl_6_n;
wire [14:0] tdl_7_n;
wire [14:0] tdl_8_n;
wire [14:0] tdl_9_n;
wire [14:0] tdl_10_n;
wire [14:0] tdl_11_n;
wire [14:0] tdl_12_n;
wire [14:0] tdl_13_n;
wire [14:0] tdl_14_n;
wire [14:0] tdl_15_n;
wire [14:0] tdl_16_n;
wire [14:0] tdl_17_n;
wire [14:0] tdl_18_n;
wire [14:0] tdl_19_n;
wire [14:0] tdl_20_n;
wire [14:0] tdl_21_n;
wire [14:0] tdl_22_n;
wire [14:0] tdl_23_n;
wire [14:0] tdl_24_n;
wire [14:0] tdl_25_n;
wire [14:0] tdl_26_n;
wire [14:0] tdl_27_n;
wire [14:0] tdl_28_n;
wire [14:0] tdl_29_n;
wire [14:0] tdl_30_n;
wire [14:0] tdl_31_n;
wire [14:0] tdl_32_n;
wire [14:0] tdl_33_n;
wire [14:0] tdl_34_n;
wire [14:0] tdl_35_n;
wire [14:0] tdl_36_n;
wire [14:0] tdl_37_n;
wire [14:0] tdl_38_n;
wire [14:0] tdl_39_n;
wire [14:0] tdl_40_n;
wire [14:0] tdl_41_n;
wire [14:0] tdl_42_n;
wire [14:0] tdl_43_n;
wire [14:0] tdl_44_n;
wire [14:0] tdl_45_n;
wire [14:0] tdl_46_n;
wire [14:0] tdl_47_n;
wire [14:0] tdl_48_n;
wire [14:0] tdl_49_n;
wire [14:0] tdl_50_n;
wire [14:0] tdl_51_n;
wire [14:0] tdl_52_n;
wire [14:0] tdl_53_n;
wire [14:0] tdl_54_n;
wire [14:0] tdl_55_n;
wire [14:0] tdl_56_n;
wire [14:0] tdl_57_n;
wire [14:0] tdl_58_n;
wire [14:0] tdl_59_n;
wire [14:0] tdl_60_n;
wire [14:0] tdl_61_n;
wire [14:0] tdl_62_n;
wire [14:0] tdl_63_n;
wire [14:0] tdl_64_n;
wire [14:0] tdl_65_n;
wire [14:0] tdl_66_n;
wire [14:0] tdl_67_n;
wire [14:0] tdl_68_n;
wire [14:0] tdl_69_n;
wire [14:0] tdl_70_n;
wire [14:0] tdl_71_n;
wire [14:0] tdl_72_n;
wire [14:0] tdl_73_n;
wire [14:0] tdl_74_n;
wire [14:0] tdl_75_n;
wire [14:0] tdl_76_n;
wire [14:0] tdl_77_n;
wire [14:0] tdl_78_n;
wire [14:0] tdl_79_n;
wire [14:0] tdl_80_n;
tdl_da_lc Utdldalc0n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(data_in), .data_out(tdl_0_n) );
defparam Utdldalc0n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc1n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_0_n), .data_out(tdl_1_n) );
defparam Utdldalc1n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc2n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_1_n), .data_out(tdl_2_n) );
defparam Utdldalc2n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc3n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_2_n), .data_out(tdl_3_n) );
defparam Utdldalc3n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc4n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_3_n), .data_out(tdl_4_n) );
defparam Utdldalc4n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc5n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_4_n), .data_out(tdl_5_n) );
defparam Utdldalc5n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc6n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_5_n), .data_out(tdl_6_n) );
defparam Utdldalc6n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc7n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_6_n), .data_out(tdl_7_n) );
defparam Utdldalc7n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc8n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_7_n), .data_out(tdl_8_n) );
defparam Utdldalc8n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc9n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_8_n), .data_out(tdl_9_n) );
defparam Utdldalc9n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc10n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_9_n), .data_out(tdl_10_n) );
defparam Utdldalc10n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc11n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_10_n), .data_out(tdl_11_n) );
defparam Utdldalc11n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc12n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_11_n), .data_out(tdl_12_n) );
defparam Utdldalc12n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc13n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_12_n), .data_out(tdl_13_n) );
defparam Utdldalc13n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc14n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_13_n), .data_out(tdl_14_n) );
defparam Utdldalc14n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc15n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_14_n), .data_out(tdl_15_n) );
defparam Utdldalc15n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc16n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_15_n), .data_out(tdl_16_n) );
defparam Utdldalc16n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc17n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_16_n), .data_out(tdl_17_n) );
defparam Utdldalc17n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc18n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_17_n), .data_out(tdl_18_n) );
defparam Utdldalc18n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc19n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_18_n), .data_out(tdl_19_n) );
defparam Utdldalc19n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc20n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_19_n), .data_out(tdl_20_n) );
defparam Utdldalc20n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc21n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_20_n), .data_out(tdl_21_n) );
defparam Utdldalc21n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc22n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_21_n), .data_out(tdl_22_n) );
defparam Utdldalc22n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc23n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_22_n), .data_out(tdl_23_n) );
defparam Utdldalc23n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc24n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_23_n), .data_out(tdl_24_n) );
defparam Utdldalc24n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc25n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_24_n), .data_out(tdl_25_n) );
defparam Utdldalc25n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc26n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_25_n), .data_out(tdl_26_n) );
defparam Utdldalc26n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc27n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_26_n), .data_out(tdl_27_n) );
defparam Utdldalc27n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc28n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_27_n), .data_out(tdl_28_n) );
defparam Utdldalc28n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc29n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_28_n), .data_out(tdl_29_n) );
defparam Utdldalc29n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc30n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_29_n), .data_out(tdl_30_n) );
defparam Utdldalc30n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc31n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_30_n), .data_out(tdl_31_n) );
defparam Utdldalc31n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc32n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_31_n), .data_out(tdl_32_n) );
defparam Utdldalc32n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc33n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_32_n), .data_out(tdl_33_n) );
defparam Utdldalc33n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc34n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_33_n), .data_out(tdl_34_n) );
defparam Utdldalc34n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc35n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_34_n), .data_out(tdl_35_n) );
defparam Utdldalc35n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc36n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_35_n), .data_out(tdl_36_n) );
defparam Utdldalc36n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc37n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_36_n), .data_out(tdl_37_n) );
defparam Utdldalc37n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc38n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_37_n), .data_out(tdl_38_n) );
defparam Utdldalc38n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc39n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_38_n), .data_out(tdl_39_n) );
defparam Utdldalc39n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc40n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_39_n), .data_out(tdl_40_n) );
defparam Utdldalc40n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc41n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_40_n), .data_out(tdl_41_n) );
defparam Utdldalc41n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc42n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_41_n), .data_out(tdl_42_n) );
defparam Utdldalc42n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc43n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_42_n), .data_out(tdl_43_n) );
defparam Utdldalc43n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc44n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_43_n), .data_out(tdl_44_n) );
defparam Utdldalc44n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc45n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_44_n), .data_out(tdl_45_n) );
defparam Utdldalc45n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc46n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_45_n), .data_out(tdl_46_n) );
defparam Utdldalc46n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc47n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_46_n), .data_out(tdl_47_n) );
defparam Utdldalc47n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc48n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_47_n), .data_out(tdl_48_n) );
defparam Utdldalc48n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc49n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_48_n), .data_out(tdl_49_n) );
defparam Utdldalc49n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc50n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_49_n), .data_out(tdl_50_n) );
defparam Utdldalc50n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc51n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_50_n), .data_out(tdl_51_n) );
defparam Utdldalc51n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc52n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_51_n), .data_out(tdl_52_n) );
defparam Utdldalc52n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc53n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_52_n), .data_out(tdl_53_n) );
defparam Utdldalc53n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc54n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_53_n), .data_out(tdl_54_n) );
defparam Utdldalc54n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc55n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_54_n), .data_out(tdl_55_n) );
defparam Utdldalc55n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc56n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_55_n), .data_out(tdl_56_n) );
defparam Utdldalc56n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc57n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_56_n), .data_out(tdl_57_n) );
defparam Utdldalc57n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc58n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_57_n), .data_out(tdl_58_n) );
defparam Utdldalc58n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc59n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_58_n), .data_out(tdl_59_n) );
defparam Utdldalc59n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc60n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_59_n), .data_out(tdl_60_n) );
defparam Utdldalc60n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc61n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_60_n), .data_out(tdl_61_n) );
defparam Utdldalc61n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc62n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_61_n), .data_out(tdl_62_n) );
defparam Utdldalc62n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc63n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_62_n), .data_out(tdl_63_n) );
defparam Utdldalc63n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc64n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_63_n), .data_out(tdl_64_n) );
defparam Utdldalc64n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc65n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_64_n), .data_out(tdl_65_n) );
defparam Utdldalc65n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc66n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_65_n), .data_out(tdl_66_n) );
defparam Utdldalc66n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc67n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_66_n), .data_out(tdl_67_n) );
defparam Utdldalc67n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc68n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_67_n), .data_out(tdl_68_n) );
defparam Utdldalc68n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc69n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_68_n), .data_out(tdl_69_n) );
defparam Utdldalc69n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc70n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_69_n), .data_out(tdl_70_n) );
defparam Utdldalc70n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc71n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_70_n), .data_out(tdl_71_n) );
defparam Utdldalc71n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc72n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_71_n), .data_out(tdl_72_n) );
defparam Utdldalc72n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc73n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_72_n), .data_out(tdl_73_n) );
defparam Utdldalc73n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc74n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_73_n), .data_out(tdl_74_n) );
defparam Utdldalc74n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc75n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_74_n), .data_out(tdl_75_n) );
defparam Utdldalc75n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc76n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_75_n), .data_out(tdl_76_n) );
defparam Utdldalc76n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc77n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_76_n), .data_out(tdl_77_n) );
defparam Utdldalc77n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc78n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_77_n), .data_out(tdl_78_n) );
defparam Utdldalc78n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc79n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_78_n), .data_out(tdl_79_n) );
defparam Utdldalc79n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc80n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_79_n), .data_out(tdl_80_n) );
defparam Utdldalc80n.WIDTH = DATA_WIDTH;
// symmetrical adders ...
wire [15:0] sym_res_0_n;
uadd_cen U_0_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_0_n), .bin(tdl_80_n), .res(sym_res_0_n) );
defparam U_0_sym_add.IN_WIDTH = 15;
defparam U_0_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_1_n;
uadd_cen U_1_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_1_n), .bin(tdl_79_n), .res(sym_res_1_n) );
defparam U_1_sym_add.IN_WIDTH = 15;
defparam U_1_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_2_n;
uadd_cen U_2_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_2_n), .bin(tdl_78_n), .res(sym_res_2_n) );
defparam U_2_sym_add.IN_WIDTH = 15;
defparam U_2_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_3_n;
uadd_cen U_3_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_3_n), .bin(tdl_77_n), .res(sym_res_3_n) );
defparam U_3_sym_add.IN_WIDTH = 15;
defparam U_3_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_4_n;
uadd_cen U_4_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_4_n), .bin(tdl_76_n), .res(sym_res_4_n) );
defparam U_4_sym_add.IN_WIDTH = 15;
defparam U_4_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_5_n;
uadd_cen U_5_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_5_n), .bin(tdl_75_n), .res(sym_res_5_n) );
defparam U_5_sym_add.IN_WIDTH = 15;
defparam U_5_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_6_n;
uadd_cen U_6_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_6_n), .bin(tdl_74_n), .res(sym_res_6_n) );
defparam U_6_sym_add.IN_WIDTH = 15;
defparam U_6_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_7_n;
uadd_cen U_7_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_7_n), .bin(tdl_73_n), .res(sym_res_7_n) );
defparam U_7_sym_add.IN_WIDTH = 15;
defparam U_7_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_8_n;
uadd_cen U_8_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_8_n), .bin(tdl_72_n), .res(sym_res_8_n) );
defparam U_8_sym_add.IN_WIDTH = 15;
defparam U_8_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_9_n;
uadd_cen U_9_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_9_n), .bin(tdl_71_n), .res(sym_res_9_n) );
defparam U_9_sym_add.IN_WIDTH = 15;
defparam U_9_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_10_n;
uadd_cen U_10_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_10_n), .bin(tdl_70_n), .res(sym_res_10_n) );
defparam U_10_sym_add.IN_WIDTH = 15;
defparam U_10_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_11_n;
uadd_cen U_11_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_11_n), .bin(tdl_69_n), .res(sym_res_11_n) );
defparam U_11_sym_add.IN_WIDTH = 15;
defparam U_11_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_12_n;
uadd_cen U_12_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_12_n), .bin(tdl_68_n), .res(sym_res_12_n) );
defparam U_12_sym_add.IN_WIDTH = 15;
defparam U_12_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_13_n;
uadd_cen U_13_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_13_n), .bin(tdl_67_n), .res(sym_res_13_n) );
defparam U_13_sym_add.IN_WIDTH = 15;
defparam U_13_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_14_n;
uadd_cen U_14_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_14_n), .bin(tdl_66_n), .res(sym_res_14_n) );
defparam U_14_sym_add.IN_WIDTH = 15;
defparam U_14_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_15_n;
uadd_cen U_15_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_15_n), .bin(tdl_65_n), .res(sym_res_15_n) );
defparam U_15_sym_add.IN_WIDTH = 15;
defparam U_15_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_16_n;
uadd_cen U_16_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_16_n), .bin(tdl_64_n), .res(sym_res_16_n) );
defparam U_16_sym_add.IN_WIDTH = 15;
defparam U_16_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_17_n;
uadd_cen U_17_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_17_n), .bin(tdl_63_n), .res(sym_res_17_n) );
defparam U_17_sym_add.IN_WIDTH = 15;
defparam U_17_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_18_n;
uadd_cen U_18_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_18_n), .bin(tdl_62_n), .res(sym_res_18_n) );
defparam U_18_sym_add.IN_WIDTH = 15;
defparam U_18_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_19_n;
uadd_cen U_19_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_19_n), .bin(tdl_61_n), .res(sym_res_19_n) );
defparam U_19_sym_add.IN_WIDTH = 15;
defparam U_19_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_20_n;
uadd_cen U_20_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_20_n), .bin(tdl_60_n), .res(sym_res_20_n) );
defparam U_20_sym_add.IN_WIDTH = 15;
defparam U_20_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_21_n;
uadd_cen U_21_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_21_n), .bin(tdl_59_n), .res(sym_res_21_n) );
defparam U_21_sym_add.IN_WIDTH = 15;
defparam U_21_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_22_n;
uadd_cen U_22_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_22_n), .bin(tdl_58_n), .res(sym_res_22_n) );
defparam U_22_sym_add.IN_WIDTH = 15;
defparam U_22_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_23_n;
uadd_cen U_23_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_23_n), .bin(tdl_57_n), .res(sym_res_23_n) );
defparam U_23_sym_add.IN_WIDTH = 15;
defparam U_23_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_24_n;
uadd_cen U_24_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_24_n), .bin(tdl_56_n), .res(sym_res_24_n) );
defparam U_24_sym_add.IN_WIDTH = 15;
defparam U_24_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_25_n;
uadd_cen U_25_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_25_n), .bin(tdl_55_n), .res(sym_res_25_n) );
defparam U_25_sym_add.IN_WIDTH = 15;
defparam U_25_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_26_n;
uadd_cen U_26_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_26_n), .bin(tdl_54_n), .res(sym_res_26_n) );
defparam U_26_sym_add.IN_WIDTH = 15;
defparam U_26_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_27_n;
uadd_cen U_27_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_27_n), .bin(tdl_53_n), .res(sym_res_27_n) );
defparam U_27_sym_add.IN_WIDTH = 15;
defparam U_27_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_28_n;
uadd_cen U_28_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_28_n), .bin(tdl_52_n), .res(sym_res_28_n) );
defparam U_28_sym_add.IN_WIDTH = 15;
defparam U_28_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_29_n;
uadd_cen U_29_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_29_n), .bin(tdl_51_n), .res(sym_res_29_n) );
defparam U_29_sym_add.IN_WIDTH = 15;
defparam U_29_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_30_n;
uadd_cen U_30_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_30_n), .bin(tdl_50_n), .res(sym_res_30_n) );
defparam U_30_sym_add.IN_WIDTH = 15;
defparam U_30_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_31_n;
uadd_cen U_31_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_31_n), .bin(tdl_49_n), .res(sym_res_31_n) );
defparam U_31_sym_add.IN_WIDTH = 15;
defparam U_31_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_32_n;
uadd_cen U_32_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_32_n), .bin(tdl_48_n), .res(sym_res_32_n) );
defparam U_32_sym_add.IN_WIDTH = 15;
defparam U_32_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_33_n;
uadd_cen U_33_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_33_n), .bin(tdl_47_n), .res(sym_res_33_n) );
defparam U_33_sym_add.IN_WIDTH = 15;
defparam U_33_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_34_n;
uadd_cen U_34_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_34_n), .bin(tdl_46_n), .res(sym_res_34_n) );
defparam U_34_sym_add.IN_WIDTH = 15;
defparam U_34_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_35_n;
uadd_cen U_35_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_35_n), .bin(tdl_45_n), .res(sym_res_35_n) );
defparam U_35_sym_add.IN_WIDTH = 15;
defparam U_35_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_36_n;
uadd_cen U_36_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_36_n), .bin(tdl_44_n), .res(sym_res_36_n) );
defparam U_36_sym_add.IN_WIDTH = 15;
defparam U_36_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_37_n;
uadd_cen U_37_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_37_n), .bin(tdl_43_n), .res(sym_res_37_n) );
defparam U_37_sym_add.IN_WIDTH = 15;
defparam U_37_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_38_n;
uadd_cen U_38_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_38_n), .bin(tdl_42_n), .res(sym_res_38_n) );
defparam U_38_sym_add.IN_WIDTH = 15;
defparam U_38_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_39_n;
uadd_cen U_39_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_39_n), .bin(tdl_41_n), .res(sym_res_39_n) );
defparam U_39_sym_add.IN_WIDTH = 15;
defparam U_39_sym_add.PIPE_DEPTH = 1;
wire [15:0] sym_res_40_n;
uadd_cen U_40_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_40_n), .bin(15'd0), .res(sym_res_40_n) );
defparam U_40_sym_add.IN_WIDTH = 15;
defparam U_40_sym_add.PIPE_DEPTH = 1;
wire [13:0] lut_val_0_n_0_pp;
rom_lut_r_cen Ur0_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[0],sym_res_2_n[0],sym_res_1_n[0],sym_res_0_n[0] } ), .data_out( lut_val_0_n_0_pp[6:0]) ) ;
 defparam Ur0_n_0_pp.DATA_WIDTH = 7;
defparam Ur0_n_0_pp.C0 = 7'd                   0;
defparam Ur0_n_0_pp.C1 = 7'd                   6;
defparam Ur0_n_0_pp.C2 = 7'd                 121;
defparam Ur0_n_0_pp.C3 = 7'd                 127;
defparam Ur0_n_0_pp.C4 = 7'd                 101;
defparam Ur0_n_0_pp.C5 = 7'd                 107;
defparam Ur0_n_0_pp.C6 = 7'd                  94;
defparam Ur0_n_0_pp.C7 = 7'd                 100;
defparam Ur0_n_0_pp.C8 = 7'd                 101;
defparam Ur0_n_0_pp.C9 = 7'd                 107;
defparam Ur0_n_0_pp.CA = 7'd                  94;
defparam Ur0_n_0_pp.CB = 7'd                 100;
defparam Ur0_n_0_pp.CC = 7'd                  74;
defparam Ur0_n_0_pp.CD = 7'd                  80;
defparam Ur0_n_0_pp.CE = 7'd                  67;
defparam Ur0_n_0_pp.CF = 7'd                  73;
assign lut_val_0_n_0_pp[13] = lut_val_0_n_0_pp[6];
assign lut_val_0_n_0_pp[12] = lut_val_0_n_0_pp[6];
assign lut_val_0_n_0_pp[11] = lut_val_0_n_0_pp[6];
assign lut_val_0_n_0_pp[10] = lut_val_0_n_0_pp[6];
assign lut_val_0_n_0_pp[9] = lut_val_0_n_0_pp[6];
assign lut_val_0_n_0_pp[8] = lut_val_0_n_0_pp[6];
assign lut_val_0_n_0_pp[7] = lut_val_0_n_0_pp[6];
wire [13:0] lut_val_0_n_1_pp;
rom_lut_r_cen Ur0_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[1],sym_res_2_n[1],sym_res_1_n[1],sym_res_0_n[1] } ), .data_out( lut_val_0_n_1_pp[6:0]) ) ;
 defparam Ur0_n_1_pp.DATA_WIDTH = 7;
defparam Ur0_n_1_pp.C0 = 7'd                   0;
defparam Ur0_n_1_pp.C1 = 7'd                   6;
defparam Ur0_n_1_pp.C2 = 7'd                 121;
defparam Ur0_n_1_pp.C3 = 7'd                 127;
defparam Ur0_n_1_pp.C4 = 7'd                 101;
defparam Ur0_n_1_pp.C5 = 7'd                 107;
defparam Ur0_n_1_pp.C6 = 7'd                  94;
defparam Ur0_n_1_pp.C7 = 7'd                 100;
defparam Ur0_n_1_pp.C8 = 7'd                 101;
defparam Ur0_n_1_pp.C9 = 7'd                 107;
defparam Ur0_n_1_pp.CA = 7'd                  94;
defparam Ur0_n_1_pp.CB = 7'd                 100;
defparam Ur0_n_1_pp.CC = 7'd                  74;
defparam Ur0_n_1_pp.CD = 7'd                  80;
defparam Ur0_n_1_pp.CE = 7'd                  67;
defparam Ur0_n_1_pp.CF = 7'd                  73;
assign lut_val_0_n_1_pp[13] = lut_val_0_n_1_pp[6];
assign lut_val_0_n_1_pp[12] = lut_val_0_n_1_pp[6];
assign lut_val_0_n_1_pp[11] = lut_val_0_n_1_pp[6];
assign lut_val_0_n_1_pp[10] = lut_val_0_n_1_pp[6];
assign lut_val_0_n_1_pp[9] = lut_val_0_n_1_pp[6];
assign lut_val_0_n_1_pp[8] = lut_val_0_n_1_pp[6];
assign lut_val_0_n_1_pp[7] = lut_val_0_n_1_pp[6];
wire [13:0] lut_val_0_n_2_pp;
rom_lut_r_cen Ur0_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[2],sym_res_2_n[2],sym_res_1_n[2],sym_res_0_n[2] } ), .data_out( lut_val_0_n_2_pp[6:0]) ) ;
 defparam Ur0_n_2_pp.DATA_WIDTH = 7;
defparam Ur0_n_2_pp.C0 = 7'd                   0;
defparam Ur0_n_2_pp.C1 = 7'd                   6;
defparam Ur0_n_2_pp.C2 = 7'd                 121;
defparam Ur0_n_2_pp.C3 = 7'd                 127;
defparam Ur0_n_2_pp.C4 = 7'd                 101;
defparam Ur0_n_2_pp.C5 = 7'd                 107;
defparam Ur0_n_2_pp.C6 = 7'd                  94;
defparam Ur0_n_2_pp.C7 = 7'd                 100;
defparam Ur0_n_2_pp.C8 = 7'd                 101;
defparam Ur0_n_2_pp.C9 = 7'd                 107;
defparam Ur0_n_2_pp.CA = 7'd                  94;
defparam Ur0_n_2_pp.CB = 7'd                 100;
defparam Ur0_n_2_pp.CC = 7'd                  74;
defparam Ur0_n_2_pp.CD = 7'd                  80;
defparam Ur0_n_2_pp.CE = 7'd                  67;
defparam Ur0_n_2_pp.CF = 7'd                  73;
assign lut_val_0_n_2_pp[13] = lut_val_0_n_2_pp[6];
assign lut_val_0_n_2_pp[12] = lut_val_0_n_2_pp[6];
assign lut_val_0_n_2_pp[11] = lut_val_0_n_2_pp[6];
assign lut_val_0_n_2_pp[10] = lut_val_0_n_2_pp[6];
assign lut_val_0_n_2_pp[9] = lut_val_0_n_2_pp[6];
assign lut_val_0_n_2_pp[8] = lut_val_0_n_2_pp[6];
assign lut_val_0_n_2_pp[7] = lut_val_0_n_2_pp[6];
wire [13:0] lut_val_0_n_3_pp;
rom_lut_r_cen Ur0_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[3],sym_res_2_n[3],sym_res_1_n[3],sym_res_0_n[3] } ), .data_out( lut_val_0_n_3_pp[6:0]) ) ;
 defparam Ur0_n_3_pp.DATA_WIDTH = 7;
defparam Ur0_n_3_pp.C0 = 7'd                   0;
defparam Ur0_n_3_pp.C1 = 7'd                   6;
defparam Ur0_n_3_pp.C2 = 7'd                 121;
defparam Ur0_n_3_pp.C3 = 7'd                 127;
defparam Ur0_n_3_pp.C4 = 7'd                 101;
defparam Ur0_n_3_pp.C5 = 7'd                 107;
defparam Ur0_n_3_pp.C6 = 7'd                  94;
defparam Ur0_n_3_pp.C7 = 7'd                 100;
defparam Ur0_n_3_pp.C8 = 7'd                 101;
defparam Ur0_n_3_pp.C9 = 7'd                 107;
defparam Ur0_n_3_pp.CA = 7'd                  94;
defparam Ur0_n_3_pp.CB = 7'd                 100;
defparam Ur0_n_3_pp.CC = 7'd                  74;
defparam Ur0_n_3_pp.CD = 7'd                  80;
defparam Ur0_n_3_pp.CE = 7'd                  67;
defparam Ur0_n_3_pp.CF = 7'd                  73;
assign lut_val_0_n_3_pp[13] = lut_val_0_n_3_pp[6];
assign lut_val_0_n_3_pp[12] = lut_val_0_n_3_pp[6];
assign lut_val_0_n_3_pp[11] = lut_val_0_n_3_pp[6];
assign lut_val_0_n_3_pp[10] = lut_val_0_n_3_pp[6];
assign lut_val_0_n_3_pp[9] = lut_val_0_n_3_pp[6];
assign lut_val_0_n_3_pp[8] = lut_val_0_n_3_pp[6];
assign lut_val_0_n_3_pp[7] = lut_val_0_n_3_pp[6];
wire [13:0] lut_val_0_n_4_pp;
rom_lut_r_cen Ur0_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[4],sym_res_2_n[4],sym_res_1_n[4],sym_res_0_n[4] } ), .data_out( lut_val_0_n_4_pp[6:0]) ) ;
 defparam Ur0_n_4_pp.DATA_WIDTH = 7;
defparam Ur0_n_4_pp.C0 = 7'd                   0;
defparam Ur0_n_4_pp.C1 = 7'd                   6;
defparam Ur0_n_4_pp.C2 = 7'd                 121;
defparam Ur0_n_4_pp.C3 = 7'd                 127;
defparam Ur0_n_4_pp.C4 = 7'd                 101;
defparam Ur0_n_4_pp.C5 = 7'd                 107;
defparam Ur0_n_4_pp.C6 = 7'd                  94;
defparam Ur0_n_4_pp.C7 = 7'd                 100;
defparam Ur0_n_4_pp.C8 = 7'd                 101;
defparam Ur0_n_4_pp.C9 = 7'd                 107;
defparam Ur0_n_4_pp.CA = 7'd                  94;
defparam Ur0_n_4_pp.CB = 7'd                 100;
defparam Ur0_n_4_pp.CC = 7'd                  74;
defparam Ur0_n_4_pp.CD = 7'd                  80;
defparam Ur0_n_4_pp.CE = 7'd                  67;
defparam Ur0_n_4_pp.CF = 7'd                  73;
assign lut_val_0_n_4_pp[13] = lut_val_0_n_4_pp[6];
assign lut_val_0_n_4_pp[12] = lut_val_0_n_4_pp[6];
assign lut_val_0_n_4_pp[11] = lut_val_0_n_4_pp[6];
assign lut_val_0_n_4_pp[10] = lut_val_0_n_4_pp[6];
assign lut_val_0_n_4_pp[9] = lut_val_0_n_4_pp[6];
assign lut_val_0_n_4_pp[8] = lut_val_0_n_4_pp[6];
assign lut_val_0_n_4_pp[7] = lut_val_0_n_4_pp[6];
wire [13:0] lut_val_0_n_5_pp;
rom_lut_r_cen Ur0_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[5],sym_res_2_n[5],sym_res_1_n[5],sym_res_0_n[5] } ), .data_out( lut_val_0_n_5_pp[6:0]) ) ;
 defparam Ur0_n_5_pp.DATA_WIDTH = 7;
defparam Ur0_n_5_pp.C0 = 7'd                   0;
defparam Ur0_n_5_pp.C1 = 7'd                   6;
defparam Ur0_n_5_pp.C2 = 7'd                 121;
defparam Ur0_n_5_pp.C3 = 7'd                 127;
defparam Ur0_n_5_pp.C4 = 7'd                 101;
defparam Ur0_n_5_pp.C5 = 7'd                 107;
defparam Ur0_n_5_pp.C6 = 7'd                  94;
defparam Ur0_n_5_pp.C7 = 7'd                 100;
defparam Ur0_n_5_pp.C8 = 7'd                 101;
defparam Ur0_n_5_pp.C9 = 7'd                 107;
defparam Ur0_n_5_pp.CA = 7'd                  94;
defparam Ur0_n_5_pp.CB = 7'd                 100;
defparam Ur0_n_5_pp.CC = 7'd                  74;
defparam Ur0_n_5_pp.CD = 7'd                  80;
defparam Ur0_n_5_pp.CE = 7'd                  67;
defparam Ur0_n_5_pp.CF = 7'd                  73;
assign lut_val_0_n_5_pp[13] = lut_val_0_n_5_pp[6];
assign lut_val_0_n_5_pp[12] = lut_val_0_n_5_pp[6];
assign lut_val_0_n_5_pp[11] = lut_val_0_n_5_pp[6];
assign lut_val_0_n_5_pp[10] = lut_val_0_n_5_pp[6];
assign lut_val_0_n_5_pp[9] = lut_val_0_n_5_pp[6];
assign lut_val_0_n_5_pp[8] = lut_val_0_n_5_pp[6];
assign lut_val_0_n_5_pp[7] = lut_val_0_n_5_pp[6];
wire [13:0] lut_val_0_n_6_pp;
rom_lut_r_cen Ur0_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[6],sym_res_2_n[6],sym_res_1_n[6],sym_res_0_n[6] } ), .data_out( lut_val_0_n_6_pp[6:0]) ) ;
 defparam Ur0_n_6_pp.DATA_WIDTH = 7;
defparam Ur0_n_6_pp.C0 = 7'd                   0;
defparam Ur0_n_6_pp.C1 = 7'd                   6;
defparam Ur0_n_6_pp.C2 = 7'd                 121;
defparam Ur0_n_6_pp.C3 = 7'd                 127;
defparam Ur0_n_6_pp.C4 = 7'd                 101;
defparam Ur0_n_6_pp.C5 = 7'd                 107;
defparam Ur0_n_6_pp.C6 = 7'd                  94;
defparam Ur0_n_6_pp.C7 = 7'd                 100;
defparam Ur0_n_6_pp.C8 = 7'd                 101;
defparam Ur0_n_6_pp.C9 = 7'd                 107;
defparam Ur0_n_6_pp.CA = 7'd                  94;
defparam Ur0_n_6_pp.CB = 7'd                 100;
defparam Ur0_n_6_pp.CC = 7'd                  74;
defparam Ur0_n_6_pp.CD = 7'd                  80;
defparam Ur0_n_6_pp.CE = 7'd                  67;
defparam Ur0_n_6_pp.CF = 7'd                  73;
assign lut_val_0_n_6_pp[13] = lut_val_0_n_6_pp[6];
assign lut_val_0_n_6_pp[12] = lut_val_0_n_6_pp[6];
assign lut_val_0_n_6_pp[11] = lut_val_0_n_6_pp[6];
assign lut_val_0_n_6_pp[10] = lut_val_0_n_6_pp[6];
assign lut_val_0_n_6_pp[9] = lut_val_0_n_6_pp[6];
assign lut_val_0_n_6_pp[8] = lut_val_0_n_6_pp[6];
assign lut_val_0_n_6_pp[7] = lut_val_0_n_6_pp[6];
wire [13:0] lut_val_0_n_7_pp;
rom_lut_r_cen Ur0_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[7],sym_res_2_n[7],sym_res_1_n[7],sym_res_0_n[7] } ), .data_out( lut_val_0_n_7_pp[6:0]) ) ;
 defparam Ur0_n_7_pp.DATA_WIDTH = 7;
defparam Ur0_n_7_pp.C0 = 7'd                   0;
defparam Ur0_n_7_pp.C1 = 7'd                   6;
defparam Ur0_n_7_pp.C2 = 7'd                 121;
defparam Ur0_n_7_pp.C3 = 7'd                 127;
defparam Ur0_n_7_pp.C4 = 7'd                 101;
defparam Ur0_n_7_pp.C5 = 7'd                 107;
defparam Ur0_n_7_pp.C6 = 7'd                  94;
defparam Ur0_n_7_pp.C7 = 7'd                 100;
defparam Ur0_n_7_pp.C8 = 7'd                 101;
defparam Ur0_n_7_pp.C9 = 7'd                 107;
defparam Ur0_n_7_pp.CA = 7'd                  94;
defparam Ur0_n_7_pp.CB = 7'd                 100;
defparam Ur0_n_7_pp.CC = 7'd                  74;
defparam Ur0_n_7_pp.CD = 7'd                  80;
defparam Ur0_n_7_pp.CE = 7'd                  67;
defparam Ur0_n_7_pp.CF = 7'd                  73;
assign lut_val_0_n_7_pp[13] = lut_val_0_n_7_pp[6];
assign lut_val_0_n_7_pp[12] = lut_val_0_n_7_pp[6];
assign lut_val_0_n_7_pp[11] = lut_val_0_n_7_pp[6];
assign lut_val_0_n_7_pp[10] = lut_val_0_n_7_pp[6];
assign lut_val_0_n_7_pp[9] = lut_val_0_n_7_pp[6];
assign lut_val_0_n_7_pp[8] = lut_val_0_n_7_pp[6];
assign lut_val_0_n_7_pp[7] = lut_val_0_n_7_pp[6];
wire [13:0] lut_val_0_n_8_pp;
rom_lut_r_cen Ur0_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[8],sym_res_2_n[8],sym_res_1_n[8],sym_res_0_n[8] } ), .data_out( lut_val_0_n_8_pp[6:0]) ) ;
 defparam Ur0_n_8_pp.DATA_WIDTH = 7;
defparam Ur0_n_8_pp.C0 = 7'd                   0;
defparam Ur0_n_8_pp.C1 = 7'd                   6;
defparam Ur0_n_8_pp.C2 = 7'd                 121;
defparam Ur0_n_8_pp.C3 = 7'd                 127;
defparam Ur0_n_8_pp.C4 = 7'd                 101;
defparam Ur0_n_8_pp.C5 = 7'd                 107;
defparam Ur0_n_8_pp.C6 = 7'd                  94;
defparam Ur0_n_8_pp.C7 = 7'd                 100;
defparam Ur0_n_8_pp.C8 = 7'd                 101;
defparam Ur0_n_8_pp.C9 = 7'd                 107;
defparam Ur0_n_8_pp.CA = 7'd                  94;
defparam Ur0_n_8_pp.CB = 7'd                 100;
defparam Ur0_n_8_pp.CC = 7'd                  74;
defparam Ur0_n_8_pp.CD = 7'd                  80;
defparam Ur0_n_8_pp.CE = 7'd                  67;
defparam Ur0_n_8_pp.CF = 7'd                  73;
assign lut_val_0_n_8_pp[13] = lut_val_0_n_8_pp[6];
assign lut_val_0_n_8_pp[12] = lut_val_0_n_8_pp[6];
assign lut_val_0_n_8_pp[11] = lut_val_0_n_8_pp[6];
assign lut_val_0_n_8_pp[10] = lut_val_0_n_8_pp[6];
assign lut_val_0_n_8_pp[9] = lut_val_0_n_8_pp[6];
assign lut_val_0_n_8_pp[8] = lut_val_0_n_8_pp[6];
assign lut_val_0_n_8_pp[7] = lut_val_0_n_8_pp[6];
wire [13:0] lut_val_0_n_9_pp;
rom_lut_r_cen Ur0_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[9],sym_res_2_n[9],sym_res_1_n[9],sym_res_0_n[9] } ), .data_out( lut_val_0_n_9_pp[6:0]) ) ;
 defparam Ur0_n_9_pp.DATA_WIDTH = 7;
defparam Ur0_n_9_pp.C0 = 7'd                   0;
defparam Ur0_n_9_pp.C1 = 7'd                   6;
defparam Ur0_n_9_pp.C2 = 7'd                 121;
defparam Ur0_n_9_pp.C3 = 7'd                 127;
defparam Ur0_n_9_pp.C4 = 7'd                 101;
defparam Ur0_n_9_pp.C5 = 7'd                 107;
defparam Ur0_n_9_pp.C6 = 7'd                  94;
defparam Ur0_n_9_pp.C7 = 7'd                 100;
defparam Ur0_n_9_pp.C8 = 7'd                 101;
defparam Ur0_n_9_pp.C9 = 7'd                 107;
defparam Ur0_n_9_pp.CA = 7'd                  94;
defparam Ur0_n_9_pp.CB = 7'd                 100;
defparam Ur0_n_9_pp.CC = 7'd                  74;
defparam Ur0_n_9_pp.CD = 7'd                  80;
defparam Ur0_n_9_pp.CE = 7'd                  67;
defparam Ur0_n_9_pp.CF = 7'd                  73;
assign lut_val_0_n_9_pp[13] = lut_val_0_n_9_pp[6];
assign lut_val_0_n_9_pp[12] = lut_val_0_n_9_pp[6];
assign lut_val_0_n_9_pp[11] = lut_val_0_n_9_pp[6];
assign lut_val_0_n_9_pp[10] = lut_val_0_n_9_pp[6];
assign lut_val_0_n_9_pp[9] = lut_val_0_n_9_pp[6];
assign lut_val_0_n_9_pp[8] = lut_val_0_n_9_pp[6];
assign lut_val_0_n_9_pp[7] = lut_val_0_n_9_pp[6];
wire [13:0] lut_val_0_n_10_pp;
rom_lut_r_cen Ur0_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[10],sym_res_2_n[10],sym_res_1_n[10],sym_res_0_n[10] } ), .data_out( lut_val_0_n_10_pp[6:0]) ) ;
 defparam Ur0_n_10_pp.DATA_WIDTH = 7;
defparam Ur0_n_10_pp.C0 = 7'd                   0;
defparam Ur0_n_10_pp.C1 = 7'd                   6;
defparam Ur0_n_10_pp.C2 = 7'd                 121;
defparam Ur0_n_10_pp.C3 = 7'd                 127;
defparam Ur0_n_10_pp.C4 = 7'd                 101;
defparam Ur0_n_10_pp.C5 = 7'd                 107;
defparam Ur0_n_10_pp.C6 = 7'd                  94;
defparam Ur0_n_10_pp.C7 = 7'd                 100;
defparam Ur0_n_10_pp.C8 = 7'd                 101;
defparam Ur0_n_10_pp.C9 = 7'd                 107;
defparam Ur0_n_10_pp.CA = 7'd                  94;
defparam Ur0_n_10_pp.CB = 7'd                 100;
defparam Ur0_n_10_pp.CC = 7'd                  74;
defparam Ur0_n_10_pp.CD = 7'd                  80;
defparam Ur0_n_10_pp.CE = 7'd                  67;
defparam Ur0_n_10_pp.CF = 7'd                  73;
assign lut_val_0_n_10_pp[13] = lut_val_0_n_10_pp[6];
assign lut_val_0_n_10_pp[12] = lut_val_0_n_10_pp[6];
assign lut_val_0_n_10_pp[11] = lut_val_0_n_10_pp[6];
assign lut_val_0_n_10_pp[10] = lut_val_0_n_10_pp[6];
assign lut_val_0_n_10_pp[9] = lut_val_0_n_10_pp[6];
assign lut_val_0_n_10_pp[8] = lut_val_0_n_10_pp[6];
assign lut_val_0_n_10_pp[7] = lut_val_0_n_10_pp[6];
wire [13:0] lut_val_0_n_11_pp;
rom_lut_r_cen Ur0_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[11],sym_res_2_n[11],sym_res_1_n[11],sym_res_0_n[11] } ), .data_out( lut_val_0_n_11_pp[6:0]) ) ;
 defparam Ur0_n_11_pp.DATA_WIDTH = 7;
defparam Ur0_n_11_pp.C0 = 7'd                   0;
defparam Ur0_n_11_pp.C1 = 7'd                   6;
defparam Ur0_n_11_pp.C2 = 7'd                 121;
defparam Ur0_n_11_pp.C3 = 7'd                 127;
defparam Ur0_n_11_pp.C4 = 7'd                 101;
defparam Ur0_n_11_pp.C5 = 7'd                 107;
defparam Ur0_n_11_pp.C6 = 7'd                  94;
defparam Ur0_n_11_pp.C7 = 7'd                 100;
defparam Ur0_n_11_pp.C8 = 7'd                 101;
defparam Ur0_n_11_pp.C9 = 7'd                 107;
defparam Ur0_n_11_pp.CA = 7'd                  94;
defparam Ur0_n_11_pp.CB = 7'd                 100;
defparam Ur0_n_11_pp.CC = 7'd                  74;
defparam Ur0_n_11_pp.CD = 7'd                  80;
defparam Ur0_n_11_pp.CE = 7'd                  67;
defparam Ur0_n_11_pp.CF = 7'd                  73;
assign lut_val_0_n_11_pp[13] = lut_val_0_n_11_pp[6];
assign lut_val_0_n_11_pp[12] = lut_val_0_n_11_pp[6];
assign lut_val_0_n_11_pp[11] = lut_val_0_n_11_pp[6];
assign lut_val_0_n_11_pp[10] = lut_val_0_n_11_pp[6];
assign lut_val_0_n_11_pp[9] = lut_val_0_n_11_pp[6];
assign lut_val_0_n_11_pp[8] = lut_val_0_n_11_pp[6];
assign lut_val_0_n_11_pp[7] = lut_val_0_n_11_pp[6];
wire [13:0] lut_val_0_n_12_pp;
rom_lut_r_cen Ur0_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[12],sym_res_2_n[12],sym_res_1_n[12],sym_res_0_n[12] } ), .data_out( lut_val_0_n_12_pp[6:0]) ) ;
 defparam Ur0_n_12_pp.DATA_WIDTH = 7;
defparam Ur0_n_12_pp.C0 = 7'd                   0;
defparam Ur0_n_12_pp.C1 = 7'd                   6;
defparam Ur0_n_12_pp.C2 = 7'd                 121;
defparam Ur0_n_12_pp.C3 = 7'd                 127;
defparam Ur0_n_12_pp.C4 = 7'd                 101;
defparam Ur0_n_12_pp.C5 = 7'd                 107;
defparam Ur0_n_12_pp.C6 = 7'd                  94;
defparam Ur0_n_12_pp.C7 = 7'd                 100;
defparam Ur0_n_12_pp.C8 = 7'd                 101;
defparam Ur0_n_12_pp.C9 = 7'd                 107;
defparam Ur0_n_12_pp.CA = 7'd                  94;
defparam Ur0_n_12_pp.CB = 7'd                 100;
defparam Ur0_n_12_pp.CC = 7'd                  74;
defparam Ur0_n_12_pp.CD = 7'd                  80;
defparam Ur0_n_12_pp.CE = 7'd                  67;
defparam Ur0_n_12_pp.CF = 7'd                  73;
assign lut_val_0_n_12_pp[13] = lut_val_0_n_12_pp[6];
assign lut_val_0_n_12_pp[12] = lut_val_0_n_12_pp[6];
assign lut_val_0_n_12_pp[11] = lut_val_0_n_12_pp[6];
assign lut_val_0_n_12_pp[10] = lut_val_0_n_12_pp[6];
assign lut_val_0_n_12_pp[9] = lut_val_0_n_12_pp[6];
assign lut_val_0_n_12_pp[8] = lut_val_0_n_12_pp[6];
assign lut_val_0_n_12_pp[7] = lut_val_0_n_12_pp[6];
wire [13:0] lut_val_0_n_13_pp;
rom_lut_r_cen Ur0_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[13],sym_res_2_n[13],sym_res_1_n[13],sym_res_0_n[13] } ), .data_out( lut_val_0_n_13_pp[6:0]) ) ;
 defparam Ur0_n_13_pp.DATA_WIDTH = 7;
defparam Ur0_n_13_pp.C0 = 7'd                   0;
defparam Ur0_n_13_pp.C1 = 7'd                   6;
defparam Ur0_n_13_pp.C2 = 7'd                 121;
defparam Ur0_n_13_pp.C3 = 7'd                 127;
defparam Ur0_n_13_pp.C4 = 7'd                 101;
defparam Ur0_n_13_pp.C5 = 7'd                 107;
defparam Ur0_n_13_pp.C6 = 7'd                  94;
defparam Ur0_n_13_pp.C7 = 7'd                 100;
defparam Ur0_n_13_pp.C8 = 7'd                 101;
defparam Ur0_n_13_pp.C9 = 7'd                 107;
defparam Ur0_n_13_pp.CA = 7'd                  94;
defparam Ur0_n_13_pp.CB = 7'd                 100;
defparam Ur0_n_13_pp.CC = 7'd                  74;
defparam Ur0_n_13_pp.CD = 7'd                  80;
defparam Ur0_n_13_pp.CE = 7'd                  67;
defparam Ur0_n_13_pp.CF = 7'd                  73;
assign lut_val_0_n_13_pp[13] = lut_val_0_n_13_pp[6];
assign lut_val_0_n_13_pp[12] = lut_val_0_n_13_pp[6];
assign lut_val_0_n_13_pp[11] = lut_val_0_n_13_pp[6];
assign lut_val_0_n_13_pp[10] = lut_val_0_n_13_pp[6];
assign lut_val_0_n_13_pp[9] = lut_val_0_n_13_pp[6];
assign lut_val_0_n_13_pp[8] = lut_val_0_n_13_pp[6];
assign lut_val_0_n_13_pp[7] = lut_val_0_n_13_pp[6];
wire [13:0] lut_val_0_n_14_pp;
rom_lut_r_cen Ur0_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[14],sym_res_2_n[14],sym_res_1_n[14],sym_res_0_n[14] } ), .data_out( lut_val_0_n_14_pp[6:0]) ) ;
 defparam Ur0_n_14_pp.DATA_WIDTH = 7;
defparam Ur0_n_14_pp.C0 = 7'd                   0;
defparam Ur0_n_14_pp.C1 = 7'd                   6;
defparam Ur0_n_14_pp.C2 = 7'd                 121;
defparam Ur0_n_14_pp.C3 = 7'd                 127;
defparam Ur0_n_14_pp.C4 = 7'd                 101;
defparam Ur0_n_14_pp.C5 = 7'd                 107;
defparam Ur0_n_14_pp.C6 = 7'd                  94;
defparam Ur0_n_14_pp.C7 = 7'd                 100;
defparam Ur0_n_14_pp.C8 = 7'd                 101;
defparam Ur0_n_14_pp.C9 = 7'd                 107;
defparam Ur0_n_14_pp.CA = 7'd                  94;
defparam Ur0_n_14_pp.CB = 7'd                 100;
defparam Ur0_n_14_pp.CC = 7'd                  74;
defparam Ur0_n_14_pp.CD = 7'd                  80;
defparam Ur0_n_14_pp.CE = 7'd                  67;
defparam Ur0_n_14_pp.CF = 7'd                  73;
assign lut_val_0_n_14_pp[13] = lut_val_0_n_14_pp[6];
assign lut_val_0_n_14_pp[12] = lut_val_0_n_14_pp[6];
assign lut_val_0_n_14_pp[11] = lut_val_0_n_14_pp[6];
assign lut_val_0_n_14_pp[10] = lut_val_0_n_14_pp[6];
assign lut_val_0_n_14_pp[9] = lut_val_0_n_14_pp[6];
assign lut_val_0_n_14_pp[8] = lut_val_0_n_14_pp[6];
assign lut_val_0_n_14_pp[7] = lut_val_0_n_14_pp[6];
wire [13:0] lut_val_0_n_15_pp;
rom_lut_r_cen Ur0_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_3_n[15],sym_res_2_n[15],sym_res_1_n[15],sym_res_0_n[15] } ), .data_out( lut_val_0_n_15_pp[6:0]) ) ;
 defparam Ur0_n_15_pp.DATA_WIDTH = 7;
defparam Ur0_n_15_pp.C0 = 7'd                   0;
defparam Ur0_n_15_pp.C1 = 7'd                   6;
defparam Ur0_n_15_pp.C2 = 7'd                 121;
defparam Ur0_n_15_pp.C3 = 7'd                 127;
defparam Ur0_n_15_pp.C4 = 7'd                 101;
defparam Ur0_n_15_pp.C5 = 7'd                 107;
defparam Ur0_n_15_pp.C6 = 7'd                  94;
defparam Ur0_n_15_pp.C7 = 7'd                 100;
defparam Ur0_n_15_pp.C8 = 7'd                 101;
defparam Ur0_n_15_pp.C9 = 7'd                 107;
defparam Ur0_n_15_pp.CA = 7'd                  94;
defparam Ur0_n_15_pp.CB = 7'd                 100;
defparam Ur0_n_15_pp.CC = 7'd                  74;
defparam Ur0_n_15_pp.CD = 7'd                  80;
defparam Ur0_n_15_pp.CE = 7'd                  67;
defparam Ur0_n_15_pp.CF = 7'd                  73;
assign lut_val_0_n_15_pp[13] = lut_val_0_n_15_pp[6];
assign lut_val_0_n_15_pp[12] = lut_val_0_n_15_pp[6];
assign lut_val_0_n_15_pp[11] = lut_val_0_n_15_pp[6];
assign lut_val_0_n_15_pp[10] = lut_val_0_n_15_pp[6];
assign lut_val_0_n_15_pp[9] = lut_val_0_n_15_pp[6];
assign lut_val_0_n_15_pp[8] = lut_val_0_n_15_pp[6];
assign lut_val_0_n_15_pp[7] = lut_val_0_n_15_pp[6];
wire [13:0] lut_val_1_n_0_pp;
rom_lut_r_cen Ur1_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[0],sym_res_6_n[0],sym_res_5_n[0],sym_res_4_n[0] } ), .data_out( lut_val_1_n_0_pp[5:0]) ) ;
 defparam Ur1_n_0_pp.DATA_WIDTH = 6;
defparam Ur1_n_0_pp.C0 = 6'd                   0;
defparam Ur1_n_0_pp.C1 = 6'd                  49;
defparam Ur1_n_0_pp.C2 = 6'd                   9;
defparam Ur1_n_0_pp.C3 = 6'd                  58;
defparam Ur1_n_0_pp.C4 = 6'd                  10;
defparam Ur1_n_0_pp.C5 = 6'd                  59;
defparam Ur1_n_0_pp.C6 = 6'd                  19;
defparam Ur1_n_0_pp.C7 = 6'd                   4;
defparam Ur1_n_0_pp.C8 = 6'd                  57;
defparam Ur1_n_0_pp.C9 = 6'd                  42;
defparam Ur1_n_0_pp.CA = 6'd                   2;
defparam Ur1_n_0_pp.CB = 6'd                  51;
defparam Ur1_n_0_pp.CC = 6'd                   3;
defparam Ur1_n_0_pp.CD = 6'd                  52;
defparam Ur1_n_0_pp.CE = 6'd                  12;
defparam Ur1_n_0_pp.CF = 6'd                  61;
assign lut_val_1_n_0_pp[13] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[12] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[11] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[10] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[9] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[8] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[7] = lut_val_1_n_0_pp[5];
assign lut_val_1_n_0_pp[6] = lut_val_1_n_0_pp[5];
wire [13:0] lut_val_1_n_1_pp;
rom_lut_r_cen Ur1_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[1],sym_res_6_n[1],sym_res_5_n[1],sym_res_4_n[1] } ), .data_out( lut_val_1_n_1_pp[5:0]) ) ;
 defparam Ur1_n_1_pp.DATA_WIDTH = 6;
defparam Ur1_n_1_pp.C0 = 6'd                   0;
defparam Ur1_n_1_pp.C1 = 6'd                  49;
defparam Ur1_n_1_pp.C2 = 6'd                   9;
defparam Ur1_n_1_pp.C3 = 6'd                  58;
defparam Ur1_n_1_pp.C4 = 6'd                  10;
defparam Ur1_n_1_pp.C5 = 6'd                  59;
defparam Ur1_n_1_pp.C6 = 6'd                  19;
defparam Ur1_n_1_pp.C7 = 6'd                   4;
defparam Ur1_n_1_pp.C8 = 6'd                  57;
defparam Ur1_n_1_pp.C9 = 6'd                  42;
defparam Ur1_n_1_pp.CA = 6'd                   2;
defparam Ur1_n_1_pp.CB = 6'd                  51;
defparam Ur1_n_1_pp.CC = 6'd                   3;
defparam Ur1_n_1_pp.CD = 6'd                  52;
defparam Ur1_n_1_pp.CE = 6'd                  12;
defparam Ur1_n_1_pp.CF = 6'd                  61;
assign lut_val_1_n_1_pp[13] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[12] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[11] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[10] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[9] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[8] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[7] = lut_val_1_n_1_pp[5];
assign lut_val_1_n_1_pp[6] = lut_val_1_n_1_pp[5];
wire [13:0] lut_val_1_n_2_pp;
rom_lut_r_cen Ur1_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[2],sym_res_6_n[2],sym_res_5_n[2],sym_res_4_n[2] } ), .data_out( lut_val_1_n_2_pp[5:0]) ) ;
 defparam Ur1_n_2_pp.DATA_WIDTH = 6;
defparam Ur1_n_2_pp.C0 = 6'd                   0;
defparam Ur1_n_2_pp.C1 = 6'd                  49;
defparam Ur1_n_2_pp.C2 = 6'd                   9;
defparam Ur1_n_2_pp.C3 = 6'd                  58;
defparam Ur1_n_2_pp.C4 = 6'd                  10;
defparam Ur1_n_2_pp.C5 = 6'd                  59;
defparam Ur1_n_2_pp.C6 = 6'd                  19;
defparam Ur1_n_2_pp.C7 = 6'd                   4;
defparam Ur1_n_2_pp.C8 = 6'd                  57;
defparam Ur1_n_2_pp.C9 = 6'd                  42;
defparam Ur1_n_2_pp.CA = 6'd                   2;
defparam Ur1_n_2_pp.CB = 6'd                  51;
defparam Ur1_n_2_pp.CC = 6'd                   3;
defparam Ur1_n_2_pp.CD = 6'd                  52;
defparam Ur1_n_2_pp.CE = 6'd                  12;
defparam Ur1_n_2_pp.CF = 6'd                  61;
assign lut_val_1_n_2_pp[13] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[12] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[11] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[10] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[9] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[8] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[7] = lut_val_1_n_2_pp[5];
assign lut_val_1_n_2_pp[6] = lut_val_1_n_2_pp[5];
wire [13:0] lut_val_1_n_3_pp;
rom_lut_r_cen Ur1_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[3],sym_res_6_n[3],sym_res_5_n[3],sym_res_4_n[3] } ), .data_out( lut_val_1_n_3_pp[5:0]) ) ;
 defparam Ur1_n_3_pp.DATA_WIDTH = 6;
defparam Ur1_n_3_pp.C0 = 6'd                   0;
defparam Ur1_n_3_pp.C1 = 6'd                  49;
defparam Ur1_n_3_pp.C2 = 6'd                   9;
defparam Ur1_n_3_pp.C3 = 6'd                  58;
defparam Ur1_n_3_pp.C4 = 6'd                  10;
defparam Ur1_n_3_pp.C5 = 6'd                  59;
defparam Ur1_n_3_pp.C6 = 6'd                  19;
defparam Ur1_n_3_pp.C7 = 6'd                   4;
defparam Ur1_n_3_pp.C8 = 6'd                  57;
defparam Ur1_n_3_pp.C9 = 6'd                  42;
defparam Ur1_n_3_pp.CA = 6'd                   2;
defparam Ur1_n_3_pp.CB = 6'd                  51;
defparam Ur1_n_3_pp.CC = 6'd                   3;
defparam Ur1_n_3_pp.CD = 6'd                  52;
defparam Ur1_n_3_pp.CE = 6'd                  12;
defparam Ur1_n_3_pp.CF = 6'd                  61;
assign lut_val_1_n_3_pp[13] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[12] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[11] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[10] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[9] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[8] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[7] = lut_val_1_n_3_pp[5];
assign lut_val_1_n_3_pp[6] = lut_val_1_n_3_pp[5];
wire [13:0] lut_val_1_n_4_pp;
rom_lut_r_cen Ur1_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[4],sym_res_6_n[4],sym_res_5_n[4],sym_res_4_n[4] } ), .data_out( lut_val_1_n_4_pp[5:0]) ) ;
 defparam Ur1_n_4_pp.DATA_WIDTH = 6;
defparam Ur1_n_4_pp.C0 = 6'd                   0;
defparam Ur1_n_4_pp.C1 = 6'd                  49;
defparam Ur1_n_4_pp.C2 = 6'd                   9;
defparam Ur1_n_4_pp.C3 = 6'd                  58;
defparam Ur1_n_4_pp.C4 = 6'd                  10;
defparam Ur1_n_4_pp.C5 = 6'd                  59;
defparam Ur1_n_4_pp.C6 = 6'd                  19;
defparam Ur1_n_4_pp.C7 = 6'd                   4;
defparam Ur1_n_4_pp.C8 = 6'd                  57;
defparam Ur1_n_4_pp.C9 = 6'd                  42;
defparam Ur1_n_4_pp.CA = 6'd                   2;
defparam Ur1_n_4_pp.CB = 6'd                  51;
defparam Ur1_n_4_pp.CC = 6'd                   3;
defparam Ur1_n_4_pp.CD = 6'd                  52;
defparam Ur1_n_4_pp.CE = 6'd                  12;
defparam Ur1_n_4_pp.CF = 6'd                  61;
assign lut_val_1_n_4_pp[13] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[12] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[11] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[10] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[9] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[8] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[7] = lut_val_1_n_4_pp[5];
assign lut_val_1_n_4_pp[6] = lut_val_1_n_4_pp[5];
wire [13:0] lut_val_1_n_5_pp;
rom_lut_r_cen Ur1_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[5],sym_res_6_n[5],sym_res_5_n[5],sym_res_4_n[5] } ), .data_out( lut_val_1_n_5_pp[5:0]) ) ;
 defparam Ur1_n_5_pp.DATA_WIDTH = 6;
defparam Ur1_n_5_pp.C0 = 6'd                   0;
defparam Ur1_n_5_pp.C1 = 6'd                  49;
defparam Ur1_n_5_pp.C2 = 6'd                   9;
defparam Ur1_n_5_pp.C3 = 6'd                  58;
defparam Ur1_n_5_pp.C4 = 6'd                  10;
defparam Ur1_n_5_pp.C5 = 6'd                  59;
defparam Ur1_n_5_pp.C6 = 6'd                  19;
defparam Ur1_n_5_pp.C7 = 6'd                   4;
defparam Ur1_n_5_pp.C8 = 6'd                  57;
defparam Ur1_n_5_pp.C9 = 6'd                  42;
defparam Ur1_n_5_pp.CA = 6'd                   2;
defparam Ur1_n_5_pp.CB = 6'd                  51;
defparam Ur1_n_5_pp.CC = 6'd                   3;
defparam Ur1_n_5_pp.CD = 6'd                  52;
defparam Ur1_n_5_pp.CE = 6'd                  12;
defparam Ur1_n_5_pp.CF = 6'd                  61;
assign lut_val_1_n_5_pp[13] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[12] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[11] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[10] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[9] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[8] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[7] = lut_val_1_n_5_pp[5];
assign lut_val_1_n_5_pp[6] = lut_val_1_n_5_pp[5];
wire [13:0] lut_val_1_n_6_pp;
rom_lut_r_cen Ur1_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[6],sym_res_6_n[6],sym_res_5_n[6],sym_res_4_n[6] } ), .data_out( lut_val_1_n_6_pp[5:0]) ) ;
 defparam Ur1_n_6_pp.DATA_WIDTH = 6;
defparam Ur1_n_6_pp.C0 = 6'd                   0;
defparam Ur1_n_6_pp.C1 = 6'd                  49;
defparam Ur1_n_6_pp.C2 = 6'd                   9;
defparam Ur1_n_6_pp.C3 = 6'd                  58;
defparam Ur1_n_6_pp.C4 = 6'd                  10;
defparam Ur1_n_6_pp.C5 = 6'd                  59;
defparam Ur1_n_6_pp.C6 = 6'd                  19;
defparam Ur1_n_6_pp.C7 = 6'd                   4;
defparam Ur1_n_6_pp.C8 = 6'd                  57;
defparam Ur1_n_6_pp.C9 = 6'd                  42;
defparam Ur1_n_6_pp.CA = 6'd                   2;
defparam Ur1_n_6_pp.CB = 6'd                  51;
defparam Ur1_n_6_pp.CC = 6'd                   3;
defparam Ur1_n_6_pp.CD = 6'd                  52;
defparam Ur1_n_6_pp.CE = 6'd                  12;
defparam Ur1_n_6_pp.CF = 6'd                  61;
assign lut_val_1_n_6_pp[13] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[12] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[11] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[10] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[9] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[8] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[7] = lut_val_1_n_6_pp[5];
assign lut_val_1_n_6_pp[6] = lut_val_1_n_6_pp[5];
wire [13:0] lut_val_1_n_7_pp;
rom_lut_r_cen Ur1_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[7],sym_res_6_n[7],sym_res_5_n[7],sym_res_4_n[7] } ), .data_out( lut_val_1_n_7_pp[5:0]) ) ;
 defparam Ur1_n_7_pp.DATA_WIDTH = 6;
defparam Ur1_n_7_pp.C0 = 6'd                   0;
defparam Ur1_n_7_pp.C1 = 6'd                  49;
defparam Ur1_n_7_pp.C2 = 6'd                   9;
defparam Ur1_n_7_pp.C3 = 6'd                  58;
defparam Ur1_n_7_pp.C4 = 6'd                  10;
defparam Ur1_n_7_pp.C5 = 6'd                  59;
defparam Ur1_n_7_pp.C6 = 6'd                  19;
defparam Ur1_n_7_pp.C7 = 6'd                   4;
defparam Ur1_n_7_pp.C8 = 6'd                  57;
defparam Ur1_n_7_pp.C9 = 6'd                  42;
defparam Ur1_n_7_pp.CA = 6'd                   2;
defparam Ur1_n_7_pp.CB = 6'd                  51;
defparam Ur1_n_7_pp.CC = 6'd                   3;
defparam Ur1_n_7_pp.CD = 6'd                  52;
defparam Ur1_n_7_pp.CE = 6'd                  12;
defparam Ur1_n_7_pp.CF = 6'd                  61;
assign lut_val_1_n_7_pp[13] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[12] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[11] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[10] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[9] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[8] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[7] = lut_val_1_n_7_pp[5];
assign lut_val_1_n_7_pp[6] = lut_val_1_n_7_pp[5];
wire [13:0] lut_val_1_n_8_pp;
rom_lut_r_cen Ur1_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[8],sym_res_6_n[8],sym_res_5_n[8],sym_res_4_n[8] } ), .data_out( lut_val_1_n_8_pp[5:0]) ) ;
 defparam Ur1_n_8_pp.DATA_WIDTH = 6;
defparam Ur1_n_8_pp.C0 = 6'd                   0;
defparam Ur1_n_8_pp.C1 = 6'd                  49;
defparam Ur1_n_8_pp.C2 = 6'd                   9;
defparam Ur1_n_8_pp.C3 = 6'd                  58;
defparam Ur1_n_8_pp.C4 = 6'd                  10;
defparam Ur1_n_8_pp.C5 = 6'd                  59;
defparam Ur1_n_8_pp.C6 = 6'd                  19;
defparam Ur1_n_8_pp.C7 = 6'd                   4;
defparam Ur1_n_8_pp.C8 = 6'd                  57;
defparam Ur1_n_8_pp.C9 = 6'd                  42;
defparam Ur1_n_8_pp.CA = 6'd                   2;
defparam Ur1_n_8_pp.CB = 6'd                  51;
defparam Ur1_n_8_pp.CC = 6'd                   3;
defparam Ur1_n_8_pp.CD = 6'd                  52;
defparam Ur1_n_8_pp.CE = 6'd                  12;
defparam Ur1_n_8_pp.CF = 6'd                  61;
assign lut_val_1_n_8_pp[13] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[12] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[11] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[10] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[9] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[8] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[7] = lut_val_1_n_8_pp[5];
assign lut_val_1_n_8_pp[6] = lut_val_1_n_8_pp[5];
wire [13:0] lut_val_1_n_9_pp;
rom_lut_r_cen Ur1_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[9],sym_res_6_n[9],sym_res_5_n[9],sym_res_4_n[9] } ), .data_out( lut_val_1_n_9_pp[5:0]) ) ;
 defparam Ur1_n_9_pp.DATA_WIDTH = 6;
defparam Ur1_n_9_pp.C0 = 6'd                   0;
defparam Ur1_n_9_pp.C1 = 6'd                  49;
defparam Ur1_n_9_pp.C2 = 6'd                   9;
defparam Ur1_n_9_pp.C3 = 6'd                  58;
defparam Ur1_n_9_pp.C4 = 6'd                  10;
defparam Ur1_n_9_pp.C5 = 6'd                  59;
defparam Ur1_n_9_pp.C6 = 6'd                  19;
defparam Ur1_n_9_pp.C7 = 6'd                   4;
defparam Ur1_n_9_pp.C8 = 6'd                  57;
defparam Ur1_n_9_pp.C9 = 6'd                  42;
defparam Ur1_n_9_pp.CA = 6'd                   2;
defparam Ur1_n_9_pp.CB = 6'd                  51;
defparam Ur1_n_9_pp.CC = 6'd                   3;
defparam Ur1_n_9_pp.CD = 6'd                  52;
defparam Ur1_n_9_pp.CE = 6'd                  12;
defparam Ur1_n_9_pp.CF = 6'd                  61;
assign lut_val_1_n_9_pp[13] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[12] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[11] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[10] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[9] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[8] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[7] = lut_val_1_n_9_pp[5];
assign lut_val_1_n_9_pp[6] = lut_val_1_n_9_pp[5];
wire [13:0] lut_val_1_n_10_pp;
rom_lut_r_cen Ur1_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[10],sym_res_6_n[10],sym_res_5_n[10],sym_res_4_n[10] } ), .data_out( lut_val_1_n_10_pp[5:0]) ) ;
 defparam Ur1_n_10_pp.DATA_WIDTH = 6;
defparam Ur1_n_10_pp.C0 = 6'd                   0;
defparam Ur1_n_10_pp.C1 = 6'd                  49;
defparam Ur1_n_10_pp.C2 = 6'd                   9;
defparam Ur1_n_10_pp.C3 = 6'd                  58;
defparam Ur1_n_10_pp.C4 = 6'd                  10;
defparam Ur1_n_10_pp.C5 = 6'd                  59;
defparam Ur1_n_10_pp.C6 = 6'd                  19;
defparam Ur1_n_10_pp.C7 = 6'd                   4;
defparam Ur1_n_10_pp.C8 = 6'd                  57;
defparam Ur1_n_10_pp.C9 = 6'd                  42;
defparam Ur1_n_10_pp.CA = 6'd                   2;
defparam Ur1_n_10_pp.CB = 6'd                  51;
defparam Ur1_n_10_pp.CC = 6'd                   3;
defparam Ur1_n_10_pp.CD = 6'd                  52;
defparam Ur1_n_10_pp.CE = 6'd                  12;
defparam Ur1_n_10_pp.CF = 6'd                  61;
assign lut_val_1_n_10_pp[13] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[12] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[11] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[10] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[9] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[8] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[7] = lut_val_1_n_10_pp[5];
assign lut_val_1_n_10_pp[6] = lut_val_1_n_10_pp[5];
wire [13:0] lut_val_1_n_11_pp;
rom_lut_r_cen Ur1_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[11],sym_res_6_n[11],sym_res_5_n[11],sym_res_4_n[11] } ), .data_out( lut_val_1_n_11_pp[5:0]) ) ;
 defparam Ur1_n_11_pp.DATA_WIDTH = 6;
defparam Ur1_n_11_pp.C0 = 6'd                   0;
defparam Ur1_n_11_pp.C1 = 6'd                  49;
defparam Ur1_n_11_pp.C2 = 6'd                   9;
defparam Ur1_n_11_pp.C3 = 6'd                  58;
defparam Ur1_n_11_pp.C4 = 6'd                  10;
defparam Ur1_n_11_pp.C5 = 6'd                  59;
defparam Ur1_n_11_pp.C6 = 6'd                  19;
defparam Ur1_n_11_pp.C7 = 6'd                   4;
defparam Ur1_n_11_pp.C8 = 6'd                  57;
defparam Ur1_n_11_pp.C9 = 6'd                  42;
defparam Ur1_n_11_pp.CA = 6'd                   2;
defparam Ur1_n_11_pp.CB = 6'd                  51;
defparam Ur1_n_11_pp.CC = 6'd                   3;
defparam Ur1_n_11_pp.CD = 6'd                  52;
defparam Ur1_n_11_pp.CE = 6'd                  12;
defparam Ur1_n_11_pp.CF = 6'd                  61;
assign lut_val_1_n_11_pp[13] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[12] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[11] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[10] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[9] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[8] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[7] = lut_val_1_n_11_pp[5];
assign lut_val_1_n_11_pp[6] = lut_val_1_n_11_pp[5];
wire [13:0] lut_val_1_n_12_pp;
rom_lut_r_cen Ur1_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[12],sym_res_6_n[12],sym_res_5_n[12],sym_res_4_n[12] } ), .data_out( lut_val_1_n_12_pp[5:0]) ) ;
 defparam Ur1_n_12_pp.DATA_WIDTH = 6;
defparam Ur1_n_12_pp.C0 = 6'd                   0;
defparam Ur1_n_12_pp.C1 = 6'd                  49;
defparam Ur1_n_12_pp.C2 = 6'd                   9;
defparam Ur1_n_12_pp.C3 = 6'd                  58;
defparam Ur1_n_12_pp.C4 = 6'd                  10;
defparam Ur1_n_12_pp.C5 = 6'd                  59;
defparam Ur1_n_12_pp.C6 = 6'd                  19;
defparam Ur1_n_12_pp.C7 = 6'd                   4;
defparam Ur1_n_12_pp.C8 = 6'd                  57;
defparam Ur1_n_12_pp.C9 = 6'd                  42;
defparam Ur1_n_12_pp.CA = 6'd                   2;
defparam Ur1_n_12_pp.CB = 6'd                  51;
defparam Ur1_n_12_pp.CC = 6'd                   3;
defparam Ur1_n_12_pp.CD = 6'd                  52;
defparam Ur1_n_12_pp.CE = 6'd                  12;
defparam Ur1_n_12_pp.CF = 6'd                  61;
assign lut_val_1_n_12_pp[13] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[12] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[11] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[10] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[9] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[8] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[7] = lut_val_1_n_12_pp[5];
assign lut_val_1_n_12_pp[6] = lut_val_1_n_12_pp[5];
wire [13:0] lut_val_1_n_13_pp;
rom_lut_r_cen Ur1_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[13],sym_res_6_n[13],sym_res_5_n[13],sym_res_4_n[13] } ), .data_out( lut_val_1_n_13_pp[5:0]) ) ;
 defparam Ur1_n_13_pp.DATA_WIDTH = 6;
defparam Ur1_n_13_pp.C0 = 6'd                   0;
defparam Ur1_n_13_pp.C1 = 6'd                  49;
defparam Ur1_n_13_pp.C2 = 6'd                   9;
defparam Ur1_n_13_pp.C3 = 6'd                  58;
defparam Ur1_n_13_pp.C4 = 6'd                  10;
defparam Ur1_n_13_pp.C5 = 6'd                  59;
defparam Ur1_n_13_pp.C6 = 6'd                  19;
defparam Ur1_n_13_pp.C7 = 6'd                   4;
defparam Ur1_n_13_pp.C8 = 6'd                  57;
defparam Ur1_n_13_pp.C9 = 6'd                  42;
defparam Ur1_n_13_pp.CA = 6'd                   2;
defparam Ur1_n_13_pp.CB = 6'd                  51;
defparam Ur1_n_13_pp.CC = 6'd                   3;
defparam Ur1_n_13_pp.CD = 6'd                  52;
defparam Ur1_n_13_pp.CE = 6'd                  12;
defparam Ur1_n_13_pp.CF = 6'd                  61;
assign lut_val_1_n_13_pp[13] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[12] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[11] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[10] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[9] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[8] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[7] = lut_val_1_n_13_pp[5];
assign lut_val_1_n_13_pp[6] = lut_val_1_n_13_pp[5];
wire [13:0] lut_val_1_n_14_pp;
rom_lut_r_cen Ur1_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[14],sym_res_6_n[14],sym_res_5_n[14],sym_res_4_n[14] } ), .data_out( lut_val_1_n_14_pp[5:0]) ) ;
 defparam Ur1_n_14_pp.DATA_WIDTH = 6;
defparam Ur1_n_14_pp.C0 = 6'd                   0;
defparam Ur1_n_14_pp.C1 = 6'd                  49;
defparam Ur1_n_14_pp.C2 = 6'd                   9;
defparam Ur1_n_14_pp.C3 = 6'd                  58;
defparam Ur1_n_14_pp.C4 = 6'd                  10;
defparam Ur1_n_14_pp.C5 = 6'd                  59;
defparam Ur1_n_14_pp.C6 = 6'd                  19;
defparam Ur1_n_14_pp.C7 = 6'd                   4;
defparam Ur1_n_14_pp.C8 = 6'd                  57;
defparam Ur1_n_14_pp.C9 = 6'd                  42;
defparam Ur1_n_14_pp.CA = 6'd                   2;
defparam Ur1_n_14_pp.CB = 6'd                  51;
defparam Ur1_n_14_pp.CC = 6'd                   3;
defparam Ur1_n_14_pp.CD = 6'd                  52;
defparam Ur1_n_14_pp.CE = 6'd                  12;
defparam Ur1_n_14_pp.CF = 6'd                  61;
assign lut_val_1_n_14_pp[13] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[12] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[11] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[10] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[9] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[8] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[7] = lut_val_1_n_14_pp[5];
assign lut_val_1_n_14_pp[6] = lut_val_1_n_14_pp[5];
wire [13:0] lut_val_1_n_15_pp;
rom_lut_r_cen Ur1_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_7_n[15],sym_res_6_n[15],sym_res_5_n[15],sym_res_4_n[15] } ), .data_out( lut_val_1_n_15_pp[5:0]) ) ;
 defparam Ur1_n_15_pp.DATA_WIDTH = 6;
defparam Ur1_n_15_pp.C0 = 6'd                   0;
defparam Ur1_n_15_pp.C1 = 6'd                  49;
defparam Ur1_n_15_pp.C2 = 6'd                   9;
defparam Ur1_n_15_pp.C3 = 6'd                  58;
defparam Ur1_n_15_pp.C4 = 6'd                  10;
defparam Ur1_n_15_pp.C5 = 6'd                  59;
defparam Ur1_n_15_pp.C6 = 6'd                  19;
defparam Ur1_n_15_pp.C7 = 6'd                   4;
defparam Ur1_n_15_pp.C8 = 6'd                  57;
defparam Ur1_n_15_pp.C9 = 6'd                  42;
defparam Ur1_n_15_pp.CA = 6'd                   2;
defparam Ur1_n_15_pp.CB = 6'd                  51;
defparam Ur1_n_15_pp.CC = 6'd                   3;
defparam Ur1_n_15_pp.CD = 6'd                  52;
defparam Ur1_n_15_pp.CE = 6'd                  12;
defparam Ur1_n_15_pp.CF = 6'd                  61;
assign lut_val_1_n_15_pp[13] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[12] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[11] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[10] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[9] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[8] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[7] = lut_val_1_n_15_pp[5];
assign lut_val_1_n_15_pp[6] = lut_val_1_n_15_pp[5];
wire [13:0] lut_val_2_n_0_pp;
rom_lut_r_cen Ur2_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[0],sym_res_10_n[0],sym_res_9_n[0],sym_res_8_n[0] } ), .data_out( lut_val_2_n_0_pp[8:0]) ) ;
 defparam Ur2_n_0_pp.DATA_WIDTH = 9;
defparam Ur2_n_0_pp.C0 = 9'd                   0;
defparam Ur2_n_0_pp.C1 = 9'd                 492;
defparam Ur2_n_0_pp.C2 = 9'd                  13;
defparam Ur2_n_0_pp.C3 = 9'd                 505;
defparam Ur2_n_0_pp.C4 = 9'd                  74;
defparam Ur2_n_0_pp.C5 = 9'd                  54;
defparam Ur2_n_0_pp.C6 = 9'd                  87;
defparam Ur2_n_0_pp.C7 = 9'd                  67;
defparam Ur2_n_0_pp.C8 = 9'd                 110;
defparam Ur2_n_0_pp.C9 = 9'd                  90;
defparam Ur2_n_0_pp.CA = 9'd                 123;
defparam Ur2_n_0_pp.CB = 9'd                 103;
defparam Ur2_n_0_pp.CC = 9'd                 184;
defparam Ur2_n_0_pp.CD = 9'd                 164;
defparam Ur2_n_0_pp.CE = 9'd                 197;
defparam Ur2_n_0_pp.CF = 9'd                 177;
assign lut_val_2_n_0_pp[13] = lut_val_2_n_0_pp[8];
assign lut_val_2_n_0_pp[12] = lut_val_2_n_0_pp[8];
assign lut_val_2_n_0_pp[11] = lut_val_2_n_0_pp[8];
assign lut_val_2_n_0_pp[10] = lut_val_2_n_0_pp[8];
assign lut_val_2_n_0_pp[9] = lut_val_2_n_0_pp[8];
wire [13:0] lut_val_2_n_1_pp;
rom_lut_r_cen Ur2_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[1],sym_res_10_n[1],sym_res_9_n[1],sym_res_8_n[1] } ), .data_out( lut_val_2_n_1_pp[8:0]) ) ;
 defparam Ur2_n_1_pp.DATA_WIDTH = 9;
defparam Ur2_n_1_pp.C0 = 9'd                   0;
defparam Ur2_n_1_pp.C1 = 9'd                 492;
defparam Ur2_n_1_pp.C2 = 9'd                  13;
defparam Ur2_n_1_pp.C3 = 9'd                 505;
defparam Ur2_n_1_pp.C4 = 9'd                  74;
defparam Ur2_n_1_pp.C5 = 9'd                  54;
defparam Ur2_n_1_pp.C6 = 9'd                  87;
defparam Ur2_n_1_pp.C7 = 9'd                  67;
defparam Ur2_n_1_pp.C8 = 9'd                 110;
defparam Ur2_n_1_pp.C9 = 9'd                  90;
defparam Ur2_n_1_pp.CA = 9'd                 123;
defparam Ur2_n_1_pp.CB = 9'd                 103;
defparam Ur2_n_1_pp.CC = 9'd                 184;
defparam Ur2_n_1_pp.CD = 9'd                 164;
defparam Ur2_n_1_pp.CE = 9'd                 197;
defparam Ur2_n_1_pp.CF = 9'd                 177;
assign lut_val_2_n_1_pp[13] = lut_val_2_n_1_pp[8];
assign lut_val_2_n_1_pp[12] = lut_val_2_n_1_pp[8];
assign lut_val_2_n_1_pp[11] = lut_val_2_n_1_pp[8];
assign lut_val_2_n_1_pp[10] = lut_val_2_n_1_pp[8];
assign lut_val_2_n_1_pp[9] = lut_val_2_n_1_pp[8];
wire [13:0] lut_val_2_n_2_pp;
rom_lut_r_cen Ur2_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[2],sym_res_10_n[2],sym_res_9_n[2],sym_res_8_n[2] } ), .data_out( lut_val_2_n_2_pp[8:0]) ) ;
 defparam Ur2_n_2_pp.DATA_WIDTH = 9;
defparam Ur2_n_2_pp.C0 = 9'd                   0;
defparam Ur2_n_2_pp.C1 = 9'd                 492;
defparam Ur2_n_2_pp.C2 = 9'd                  13;
defparam Ur2_n_2_pp.C3 = 9'd                 505;
defparam Ur2_n_2_pp.C4 = 9'd                  74;
defparam Ur2_n_2_pp.C5 = 9'd                  54;
defparam Ur2_n_2_pp.C6 = 9'd                  87;
defparam Ur2_n_2_pp.C7 = 9'd                  67;
defparam Ur2_n_2_pp.C8 = 9'd                 110;
defparam Ur2_n_2_pp.C9 = 9'd                  90;
defparam Ur2_n_2_pp.CA = 9'd                 123;
defparam Ur2_n_2_pp.CB = 9'd                 103;
defparam Ur2_n_2_pp.CC = 9'd                 184;
defparam Ur2_n_2_pp.CD = 9'd                 164;
defparam Ur2_n_2_pp.CE = 9'd                 197;
defparam Ur2_n_2_pp.CF = 9'd                 177;
assign lut_val_2_n_2_pp[13] = lut_val_2_n_2_pp[8];
assign lut_val_2_n_2_pp[12] = lut_val_2_n_2_pp[8];
assign lut_val_2_n_2_pp[11] = lut_val_2_n_2_pp[8];
assign lut_val_2_n_2_pp[10] = lut_val_2_n_2_pp[8];
assign lut_val_2_n_2_pp[9] = lut_val_2_n_2_pp[8];
wire [13:0] lut_val_2_n_3_pp;
rom_lut_r_cen Ur2_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[3],sym_res_10_n[3],sym_res_9_n[3],sym_res_8_n[3] } ), .data_out( lut_val_2_n_3_pp[8:0]) ) ;
 defparam Ur2_n_3_pp.DATA_WIDTH = 9;
defparam Ur2_n_3_pp.C0 = 9'd                   0;
defparam Ur2_n_3_pp.C1 = 9'd                 492;
defparam Ur2_n_3_pp.C2 = 9'd                  13;
defparam Ur2_n_3_pp.C3 = 9'd                 505;
defparam Ur2_n_3_pp.C4 = 9'd                  74;
defparam Ur2_n_3_pp.C5 = 9'd                  54;
defparam Ur2_n_3_pp.C6 = 9'd                  87;
defparam Ur2_n_3_pp.C7 = 9'd                  67;
defparam Ur2_n_3_pp.C8 = 9'd                 110;
defparam Ur2_n_3_pp.C9 = 9'd                  90;
defparam Ur2_n_3_pp.CA = 9'd                 123;
defparam Ur2_n_3_pp.CB = 9'd                 103;
defparam Ur2_n_3_pp.CC = 9'd                 184;
defparam Ur2_n_3_pp.CD = 9'd                 164;
defparam Ur2_n_3_pp.CE = 9'd                 197;
defparam Ur2_n_3_pp.CF = 9'd                 177;
assign lut_val_2_n_3_pp[13] = lut_val_2_n_3_pp[8];
assign lut_val_2_n_3_pp[12] = lut_val_2_n_3_pp[8];
assign lut_val_2_n_3_pp[11] = lut_val_2_n_3_pp[8];
assign lut_val_2_n_3_pp[10] = lut_val_2_n_3_pp[8];
assign lut_val_2_n_3_pp[9] = lut_val_2_n_3_pp[8];
wire [13:0] lut_val_2_n_4_pp;
rom_lut_r_cen Ur2_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[4],sym_res_10_n[4],sym_res_9_n[4],sym_res_8_n[4] } ), .data_out( lut_val_2_n_4_pp[8:0]) ) ;
 defparam Ur2_n_4_pp.DATA_WIDTH = 9;
defparam Ur2_n_4_pp.C0 = 9'd                   0;
defparam Ur2_n_4_pp.C1 = 9'd                 492;
defparam Ur2_n_4_pp.C2 = 9'd                  13;
defparam Ur2_n_4_pp.C3 = 9'd                 505;
defparam Ur2_n_4_pp.C4 = 9'd                  74;
defparam Ur2_n_4_pp.C5 = 9'd                  54;
defparam Ur2_n_4_pp.C6 = 9'd                  87;
defparam Ur2_n_4_pp.C7 = 9'd                  67;
defparam Ur2_n_4_pp.C8 = 9'd                 110;
defparam Ur2_n_4_pp.C9 = 9'd                  90;
defparam Ur2_n_4_pp.CA = 9'd                 123;
defparam Ur2_n_4_pp.CB = 9'd                 103;
defparam Ur2_n_4_pp.CC = 9'd                 184;
defparam Ur2_n_4_pp.CD = 9'd                 164;
defparam Ur2_n_4_pp.CE = 9'd                 197;
defparam Ur2_n_4_pp.CF = 9'd                 177;
assign lut_val_2_n_4_pp[13] = lut_val_2_n_4_pp[8];
assign lut_val_2_n_4_pp[12] = lut_val_2_n_4_pp[8];
assign lut_val_2_n_4_pp[11] = lut_val_2_n_4_pp[8];
assign lut_val_2_n_4_pp[10] = lut_val_2_n_4_pp[8];
assign lut_val_2_n_4_pp[9] = lut_val_2_n_4_pp[8];
wire [13:0] lut_val_2_n_5_pp;
rom_lut_r_cen Ur2_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[5],sym_res_10_n[5],sym_res_9_n[5],sym_res_8_n[5] } ), .data_out( lut_val_2_n_5_pp[8:0]) ) ;
 defparam Ur2_n_5_pp.DATA_WIDTH = 9;
defparam Ur2_n_5_pp.C0 = 9'd                   0;
defparam Ur2_n_5_pp.C1 = 9'd                 492;
defparam Ur2_n_5_pp.C2 = 9'd                  13;
defparam Ur2_n_5_pp.C3 = 9'd                 505;
defparam Ur2_n_5_pp.C4 = 9'd                  74;
defparam Ur2_n_5_pp.C5 = 9'd                  54;
defparam Ur2_n_5_pp.C6 = 9'd                  87;
defparam Ur2_n_5_pp.C7 = 9'd                  67;
defparam Ur2_n_5_pp.C8 = 9'd                 110;
defparam Ur2_n_5_pp.C9 = 9'd                  90;
defparam Ur2_n_5_pp.CA = 9'd                 123;
defparam Ur2_n_5_pp.CB = 9'd                 103;
defparam Ur2_n_5_pp.CC = 9'd                 184;
defparam Ur2_n_5_pp.CD = 9'd                 164;
defparam Ur2_n_5_pp.CE = 9'd                 197;
defparam Ur2_n_5_pp.CF = 9'd                 177;
assign lut_val_2_n_5_pp[13] = lut_val_2_n_5_pp[8];
assign lut_val_2_n_5_pp[12] = lut_val_2_n_5_pp[8];
assign lut_val_2_n_5_pp[11] = lut_val_2_n_5_pp[8];
assign lut_val_2_n_5_pp[10] = lut_val_2_n_5_pp[8];
assign lut_val_2_n_5_pp[9] = lut_val_2_n_5_pp[8];
wire [13:0] lut_val_2_n_6_pp;
rom_lut_r_cen Ur2_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[6],sym_res_10_n[6],sym_res_9_n[6],sym_res_8_n[6] } ), .data_out( lut_val_2_n_6_pp[8:0]) ) ;
 defparam Ur2_n_6_pp.DATA_WIDTH = 9;
defparam Ur2_n_6_pp.C0 = 9'd                   0;
defparam Ur2_n_6_pp.C1 = 9'd                 492;
defparam Ur2_n_6_pp.C2 = 9'd                  13;
defparam Ur2_n_6_pp.C3 = 9'd                 505;
defparam Ur2_n_6_pp.C4 = 9'd                  74;
defparam Ur2_n_6_pp.C5 = 9'd                  54;
defparam Ur2_n_6_pp.C6 = 9'd                  87;
defparam Ur2_n_6_pp.C7 = 9'd                  67;
defparam Ur2_n_6_pp.C8 = 9'd                 110;
defparam Ur2_n_6_pp.C9 = 9'd                  90;
defparam Ur2_n_6_pp.CA = 9'd                 123;
defparam Ur2_n_6_pp.CB = 9'd                 103;
defparam Ur2_n_6_pp.CC = 9'd                 184;
defparam Ur2_n_6_pp.CD = 9'd                 164;
defparam Ur2_n_6_pp.CE = 9'd                 197;
defparam Ur2_n_6_pp.CF = 9'd                 177;
assign lut_val_2_n_6_pp[13] = lut_val_2_n_6_pp[8];
assign lut_val_2_n_6_pp[12] = lut_val_2_n_6_pp[8];
assign lut_val_2_n_6_pp[11] = lut_val_2_n_6_pp[8];
assign lut_val_2_n_6_pp[10] = lut_val_2_n_6_pp[8];
assign lut_val_2_n_6_pp[9] = lut_val_2_n_6_pp[8];
wire [13:0] lut_val_2_n_7_pp;
rom_lut_r_cen Ur2_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[7],sym_res_10_n[7],sym_res_9_n[7],sym_res_8_n[7] } ), .data_out( lut_val_2_n_7_pp[8:0]) ) ;
 defparam Ur2_n_7_pp.DATA_WIDTH = 9;
defparam Ur2_n_7_pp.C0 = 9'd                   0;
defparam Ur2_n_7_pp.C1 = 9'd                 492;
defparam Ur2_n_7_pp.C2 = 9'd                  13;
defparam Ur2_n_7_pp.C3 = 9'd                 505;
defparam Ur2_n_7_pp.C4 = 9'd                  74;
defparam Ur2_n_7_pp.C5 = 9'd                  54;
defparam Ur2_n_7_pp.C6 = 9'd                  87;
defparam Ur2_n_7_pp.C7 = 9'd                  67;
defparam Ur2_n_7_pp.C8 = 9'd                 110;
defparam Ur2_n_7_pp.C9 = 9'd                  90;
defparam Ur2_n_7_pp.CA = 9'd                 123;
defparam Ur2_n_7_pp.CB = 9'd                 103;
defparam Ur2_n_7_pp.CC = 9'd                 184;
defparam Ur2_n_7_pp.CD = 9'd                 164;
defparam Ur2_n_7_pp.CE = 9'd                 197;
defparam Ur2_n_7_pp.CF = 9'd                 177;
assign lut_val_2_n_7_pp[13] = lut_val_2_n_7_pp[8];
assign lut_val_2_n_7_pp[12] = lut_val_2_n_7_pp[8];
assign lut_val_2_n_7_pp[11] = lut_val_2_n_7_pp[8];
assign lut_val_2_n_7_pp[10] = lut_val_2_n_7_pp[8];
assign lut_val_2_n_7_pp[9] = lut_val_2_n_7_pp[8];
wire [13:0] lut_val_2_n_8_pp;
rom_lut_r_cen Ur2_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[8],sym_res_10_n[8],sym_res_9_n[8],sym_res_8_n[8] } ), .data_out( lut_val_2_n_8_pp[8:0]) ) ;
 defparam Ur2_n_8_pp.DATA_WIDTH = 9;
defparam Ur2_n_8_pp.C0 = 9'd                   0;
defparam Ur2_n_8_pp.C1 = 9'd                 492;
defparam Ur2_n_8_pp.C2 = 9'd                  13;
defparam Ur2_n_8_pp.C3 = 9'd                 505;
defparam Ur2_n_8_pp.C4 = 9'd                  74;
defparam Ur2_n_8_pp.C5 = 9'd                  54;
defparam Ur2_n_8_pp.C6 = 9'd                  87;
defparam Ur2_n_8_pp.C7 = 9'd                  67;
defparam Ur2_n_8_pp.C8 = 9'd                 110;
defparam Ur2_n_8_pp.C9 = 9'd                  90;
defparam Ur2_n_8_pp.CA = 9'd                 123;
defparam Ur2_n_8_pp.CB = 9'd                 103;
defparam Ur2_n_8_pp.CC = 9'd                 184;
defparam Ur2_n_8_pp.CD = 9'd                 164;
defparam Ur2_n_8_pp.CE = 9'd                 197;
defparam Ur2_n_8_pp.CF = 9'd                 177;
assign lut_val_2_n_8_pp[13] = lut_val_2_n_8_pp[8];
assign lut_val_2_n_8_pp[12] = lut_val_2_n_8_pp[8];
assign lut_val_2_n_8_pp[11] = lut_val_2_n_8_pp[8];
assign lut_val_2_n_8_pp[10] = lut_val_2_n_8_pp[8];
assign lut_val_2_n_8_pp[9] = lut_val_2_n_8_pp[8];
wire [13:0] lut_val_2_n_9_pp;
rom_lut_r_cen Ur2_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[9],sym_res_10_n[9],sym_res_9_n[9],sym_res_8_n[9] } ), .data_out( lut_val_2_n_9_pp[8:0]) ) ;
 defparam Ur2_n_9_pp.DATA_WIDTH = 9;
defparam Ur2_n_9_pp.C0 = 9'd                   0;
defparam Ur2_n_9_pp.C1 = 9'd                 492;
defparam Ur2_n_9_pp.C2 = 9'd                  13;
defparam Ur2_n_9_pp.C3 = 9'd                 505;
defparam Ur2_n_9_pp.C4 = 9'd                  74;
defparam Ur2_n_9_pp.C5 = 9'd                  54;
defparam Ur2_n_9_pp.C6 = 9'd                  87;
defparam Ur2_n_9_pp.C7 = 9'd                  67;
defparam Ur2_n_9_pp.C8 = 9'd                 110;
defparam Ur2_n_9_pp.C9 = 9'd                  90;
defparam Ur2_n_9_pp.CA = 9'd                 123;
defparam Ur2_n_9_pp.CB = 9'd                 103;
defparam Ur2_n_9_pp.CC = 9'd                 184;
defparam Ur2_n_9_pp.CD = 9'd                 164;
defparam Ur2_n_9_pp.CE = 9'd                 197;
defparam Ur2_n_9_pp.CF = 9'd                 177;
assign lut_val_2_n_9_pp[13] = lut_val_2_n_9_pp[8];
assign lut_val_2_n_9_pp[12] = lut_val_2_n_9_pp[8];
assign lut_val_2_n_9_pp[11] = lut_val_2_n_9_pp[8];
assign lut_val_2_n_9_pp[10] = lut_val_2_n_9_pp[8];
assign lut_val_2_n_9_pp[9] = lut_val_2_n_9_pp[8];
wire [13:0] lut_val_2_n_10_pp;
rom_lut_r_cen Ur2_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[10],sym_res_10_n[10],sym_res_9_n[10],sym_res_8_n[10] } ), .data_out( lut_val_2_n_10_pp[8:0]) ) ;
 defparam Ur2_n_10_pp.DATA_WIDTH = 9;
defparam Ur2_n_10_pp.C0 = 9'd                   0;
defparam Ur2_n_10_pp.C1 = 9'd                 492;
defparam Ur2_n_10_pp.C2 = 9'd                  13;
defparam Ur2_n_10_pp.C3 = 9'd                 505;
defparam Ur2_n_10_pp.C4 = 9'd                  74;
defparam Ur2_n_10_pp.C5 = 9'd                  54;
defparam Ur2_n_10_pp.C6 = 9'd                  87;
defparam Ur2_n_10_pp.C7 = 9'd                  67;
defparam Ur2_n_10_pp.C8 = 9'd                 110;
defparam Ur2_n_10_pp.C9 = 9'd                  90;
defparam Ur2_n_10_pp.CA = 9'd                 123;
defparam Ur2_n_10_pp.CB = 9'd                 103;
defparam Ur2_n_10_pp.CC = 9'd                 184;
defparam Ur2_n_10_pp.CD = 9'd                 164;
defparam Ur2_n_10_pp.CE = 9'd                 197;
defparam Ur2_n_10_pp.CF = 9'd                 177;
assign lut_val_2_n_10_pp[13] = lut_val_2_n_10_pp[8];
assign lut_val_2_n_10_pp[12] = lut_val_2_n_10_pp[8];
assign lut_val_2_n_10_pp[11] = lut_val_2_n_10_pp[8];
assign lut_val_2_n_10_pp[10] = lut_val_2_n_10_pp[8];
assign lut_val_2_n_10_pp[9] = lut_val_2_n_10_pp[8];
wire [13:0] lut_val_2_n_11_pp;
rom_lut_r_cen Ur2_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[11],sym_res_10_n[11],sym_res_9_n[11],sym_res_8_n[11] } ), .data_out( lut_val_2_n_11_pp[8:0]) ) ;
 defparam Ur2_n_11_pp.DATA_WIDTH = 9;
defparam Ur2_n_11_pp.C0 = 9'd                   0;
defparam Ur2_n_11_pp.C1 = 9'd                 492;
defparam Ur2_n_11_pp.C2 = 9'd                  13;
defparam Ur2_n_11_pp.C3 = 9'd                 505;
defparam Ur2_n_11_pp.C4 = 9'd                  74;
defparam Ur2_n_11_pp.C5 = 9'd                  54;
defparam Ur2_n_11_pp.C6 = 9'd                  87;
defparam Ur2_n_11_pp.C7 = 9'd                  67;
defparam Ur2_n_11_pp.C8 = 9'd                 110;
defparam Ur2_n_11_pp.C9 = 9'd                  90;
defparam Ur2_n_11_pp.CA = 9'd                 123;
defparam Ur2_n_11_pp.CB = 9'd                 103;
defparam Ur2_n_11_pp.CC = 9'd                 184;
defparam Ur2_n_11_pp.CD = 9'd                 164;
defparam Ur2_n_11_pp.CE = 9'd                 197;
defparam Ur2_n_11_pp.CF = 9'd                 177;
assign lut_val_2_n_11_pp[13] = lut_val_2_n_11_pp[8];
assign lut_val_2_n_11_pp[12] = lut_val_2_n_11_pp[8];
assign lut_val_2_n_11_pp[11] = lut_val_2_n_11_pp[8];
assign lut_val_2_n_11_pp[10] = lut_val_2_n_11_pp[8];
assign lut_val_2_n_11_pp[9] = lut_val_2_n_11_pp[8];
wire [13:0] lut_val_2_n_12_pp;
rom_lut_r_cen Ur2_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[12],sym_res_10_n[12],sym_res_9_n[12],sym_res_8_n[12] } ), .data_out( lut_val_2_n_12_pp[8:0]) ) ;
 defparam Ur2_n_12_pp.DATA_WIDTH = 9;
defparam Ur2_n_12_pp.C0 = 9'd                   0;
defparam Ur2_n_12_pp.C1 = 9'd                 492;
defparam Ur2_n_12_pp.C2 = 9'd                  13;
defparam Ur2_n_12_pp.C3 = 9'd                 505;
defparam Ur2_n_12_pp.C4 = 9'd                  74;
defparam Ur2_n_12_pp.C5 = 9'd                  54;
defparam Ur2_n_12_pp.C6 = 9'd                  87;
defparam Ur2_n_12_pp.C7 = 9'd                  67;
defparam Ur2_n_12_pp.C8 = 9'd                 110;
defparam Ur2_n_12_pp.C9 = 9'd                  90;
defparam Ur2_n_12_pp.CA = 9'd                 123;
defparam Ur2_n_12_pp.CB = 9'd                 103;
defparam Ur2_n_12_pp.CC = 9'd                 184;
defparam Ur2_n_12_pp.CD = 9'd                 164;
defparam Ur2_n_12_pp.CE = 9'd                 197;
defparam Ur2_n_12_pp.CF = 9'd                 177;
assign lut_val_2_n_12_pp[13] = lut_val_2_n_12_pp[8];
assign lut_val_2_n_12_pp[12] = lut_val_2_n_12_pp[8];
assign lut_val_2_n_12_pp[11] = lut_val_2_n_12_pp[8];
assign lut_val_2_n_12_pp[10] = lut_val_2_n_12_pp[8];
assign lut_val_2_n_12_pp[9] = lut_val_2_n_12_pp[8];
wire [13:0] lut_val_2_n_13_pp;
rom_lut_r_cen Ur2_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[13],sym_res_10_n[13],sym_res_9_n[13],sym_res_8_n[13] } ), .data_out( lut_val_2_n_13_pp[8:0]) ) ;
 defparam Ur2_n_13_pp.DATA_WIDTH = 9;
defparam Ur2_n_13_pp.C0 = 9'd                   0;
defparam Ur2_n_13_pp.C1 = 9'd                 492;
defparam Ur2_n_13_pp.C2 = 9'd                  13;
defparam Ur2_n_13_pp.C3 = 9'd                 505;
defparam Ur2_n_13_pp.C4 = 9'd                  74;
defparam Ur2_n_13_pp.C5 = 9'd                  54;
defparam Ur2_n_13_pp.C6 = 9'd                  87;
defparam Ur2_n_13_pp.C7 = 9'd                  67;
defparam Ur2_n_13_pp.C8 = 9'd                 110;
defparam Ur2_n_13_pp.C9 = 9'd                  90;
defparam Ur2_n_13_pp.CA = 9'd                 123;
defparam Ur2_n_13_pp.CB = 9'd                 103;
defparam Ur2_n_13_pp.CC = 9'd                 184;
defparam Ur2_n_13_pp.CD = 9'd                 164;
defparam Ur2_n_13_pp.CE = 9'd                 197;
defparam Ur2_n_13_pp.CF = 9'd                 177;
assign lut_val_2_n_13_pp[13] = lut_val_2_n_13_pp[8];
assign lut_val_2_n_13_pp[12] = lut_val_2_n_13_pp[8];
assign lut_val_2_n_13_pp[11] = lut_val_2_n_13_pp[8];
assign lut_val_2_n_13_pp[10] = lut_val_2_n_13_pp[8];
assign lut_val_2_n_13_pp[9] = lut_val_2_n_13_pp[8];
wire [13:0] lut_val_2_n_14_pp;
rom_lut_r_cen Ur2_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[14],sym_res_10_n[14],sym_res_9_n[14],sym_res_8_n[14] } ), .data_out( lut_val_2_n_14_pp[8:0]) ) ;
 defparam Ur2_n_14_pp.DATA_WIDTH = 9;
defparam Ur2_n_14_pp.C0 = 9'd                   0;
defparam Ur2_n_14_pp.C1 = 9'd                 492;
defparam Ur2_n_14_pp.C2 = 9'd                  13;
defparam Ur2_n_14_pp.C3 = 9'd                 505;
defparam Ur2_n_14_pp.C4 = 9'd                  74;
defparam Ur2_n_14_pp.C5 = 9'd                  54;
defparam Ur2_n_14_pp.C6 = 9'd                  87;
defparam Ur2_n_14_pp.C7 = 9'd                  67;
defparam Ur2_n_14_pp.C8 = 9'd                 110;
defparam Ur2_n_14_pp.C9 = 9'd                  90;
defparam Ur2_n_14_pp.CA = 9'd                 123;
defparam Ur2_n_14_pp.CB = 9'd                 103;
defparam Ur2_n_14_pp.CC = 9'd                 184;
defparam Ur2_n_14_pp.CD = 9'd                 164;
defparam Ur2_n_14_pp.CE = 9'd                 197;
defparam Ur2_n_14_pp.CF = 9'd                 177;
assign lut_val_2_n_14_pp[13] = lut_val_2_n_14_pp[8];
assign lut_val_2_n_14_pp[12] = lut_val_2_n_14_pp[8];
assign lut_val_2_n_14_pp[11] = lut_val_2_n_14_pp[8];
assign lut_val_2_n_14_pp[10] = lut_val_2_n_14_pp[8];
assign lut_val_2_n_14_pp[9] = lut_val_2_n_14_pp[8];
wire [13:0] lut_val_2_n_15_pp;
rom_lut_r_cen Ur2_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_11_n[15],sym_res_10_n[15],sym_res_9_n[15],sym_res_8_n[15] } ), .data_out( lut_val_2_n_15_pp[8:0]) ) ;
 defparam Ur2_n_15_pp.DATA_WIDTH = 9;
defparam Ur2_n_15_pp.C0 = 9'd                   0;
defparam Ur2_n_15_pp.C1 = 9'd                 492;
defparam Ur2_n_15_pp.C2 = 9'd                  13;
defparam Ur2_n_15_pp.C3 = 9'd                 505;
defparam Ur2_n_15_pp.C4 = 9'd                  74;
defparam Ur2_n_15_pp.C5 = 9'd                  54;
defparam Ur2_n_15_pp.C6 = 9'd                  87;
defparam Ur2_n_15_pp.C7 = 9'd                  67;
defparam Ur2_n_15_pp.C8 = 9'd                 110;
defparam Ur2_n_15_pp.C9 = 9'd                  90;
defparam Ur2_n_15_pp.CA = 9'd                 123;
defparam Ur2_n_15_pp.CB = 9'd                 103;
defparam Ur2_n_15_pp.CC = 9'd                 184;
defparam Ur2_n_15_pp.CD = 9'd                 164;
defparam Ur2_n_15_pp.CE = 9'd                 197;
defparam Ur2_n_15_pp.CF = 9'd                 177;
assign lut_val_2_n_15_pp[13] = lut_val_2_n_15_pp[8];
assign lut_val_2_n_15_pp[12] = lut_val_2_n_15_pp[8];
assign lut_val_2_n_15_pp[11] = lut_val_2_n_15_pp[8];
assign lut_val_2_n_15_pp[10] = lut_val_2_n_15_pp[8];
assign lut_val_2_n_15_pp[9] = lut_val_2_n_15_pp[8];
wire [13:0] lut_val_3_n_0_pp;
rom_lut_r_cen Ur3_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[0],sym_res_14_n[0],sym_res_13_n[0],sym_res_12_n[0] } ), .data_out( lut_val_3_n_0_pp[7:0]) ) ;
 defparam Ur3_n_0_pp.DATA_WIDTH = 8;
defparam Ur3_n_0_pp.C0 = 8'd                   0;
defparam Ur3_n_0_pp.C1 = 8'd                  72;
defparam Ur3_n_0_pp.C2 = 8'd                 251;
defparam Ur3_n_0_pp.C3 = 8'd                  67;
defparam Ur3_n_0_pp.C4 = 8'd                 214;
defparam Ur3_n_0_pp.C5 = 8'd                  30;
defparam Ur3_n_0_pp.C6 = 8'd                 209;
defparam Ur3_n_0_pp.C7 = 8'd                  25;
defparam Ur3_n_0_pp.C8 = 8'd                   1;
defparam Ur3_n_0_pp.C9 = 8'd                  73;
defparam Ur3_n_0_pp.CA = 8'd                 252;
defparam Ur3_n_0_pp.CB = 8'd                  68;
defparam Ur3_n_0_pp.CC = 8'd                 215;
defparam Ur3_n_0_pp.CD = 8'd                  31;
defparam Ur3_n_0_pp.CE = 8'd                 210;
defparam Ur3_n_0_pp.CF = 8'd                  26;
assign lut_val_3_n_0_pp[13] = lut_val_3_n_0_pp[7];
assign lut_val_3_n_0_pp[12] = lut_val_3_n_0_pp[7];
assign lut_val_3_n_0_pp[11] = lut_val_3_n_0_pp[7];
assign lut_val_3_n_0_pp[10] = lut_val_3_n_0_pp[7];
assign lut_val_3_n_0_pp[9] = lut_val_3_n_0_pp[7];
assign lut_val_3_n_0_pp[8] = lut_val_3_n_0_pp[7];
wire [13:0] lut_val_3_n_1_pp;
rom_lut_r_cen Ur3_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[1],sym_res_14_n[1],sym_res_13_n[1],sym_res_12_n[1] } ), .data_out( lut_val_3_n_1_pp[7:0]) ) ;
 defparam Ur3_n_1_pp.DATA_WIDTH = 8;
defparam Ur3_n_1_pp.C0 = 8'd                   0;
defparam Ur3_n_1_pp.C1 = 8'd                  72;
defparam Ur3_n_1_pp.C2 = 8'd                 251;
defparam Ur3_n_1_pp.C3 = 8'd                  67;
defparam Ur3_n_1_pp.C4 = 8'd                 214;
defparam Ur3_n_1_pp.C5 = 8'd                  30;
defparam Ur3_n_1_pp.C6 = 8'd                 209;
defparam Ur3_n_1_pp.C7 = 8'd                  25;
defparam Ur3_n_1_pp.C8 = 8'd                   1;
defparam Ur3_n_1_pp.C9 = 8'd                  73;
defparam Ur3_n_1_pp.CA = 8'd                 252;
defparam Ur3_n_1_pp.CB = 8'd                  68;
defparam Ur3_n_1_pp.CC = 8'd                 215;
defparam Ur3_n_1_pp.CD = 8'd                  31;
defparam Ur3_n_1_pp.CE = 8'd                 210;
defparam Ur3_n_1_pp.CF = 8'd                  26;
assign lut_val_3_n_1_pp[13] = lut_val_3_n_1_pp[7];
assign lut_val_3_n_1_pp[12] = lut_val_3_n_1_pp[7];
assign lut_val_3_n_1_pp[11] = lut_val_3_n_1_pp[7];
assign lut_val_3_n_1_pp[10] = lut_val_3_n_1_pp[7];
assign lut_val_3_n_1_pp[9] = lut_val_3_n_1_pp[7];
assign lut_val_3_n_1_pp[8] = lut_val_3_n_1_pp[7];
wire [13:0] lut_val_3_n_2_pp;
rom_lut_r_cen Ur3_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[2],sym_res_14_n[2],sym_res_13_n[2],sym_res_12_n[2] } ), .data_out( lut_val_3_n_2_pp[7:0]) ) ;
 defparam Ur3_n_2_pp.DATA_WIDTH = 8;
defparam Ur3_n_2_pp.C0 = 8'd                   0;
defparam Ur3_n_2_pp.C1 = 8'd                  72;
defparam Ur3_n_2_pp.C2 = 8'd                 251;
defparam Ur3_n_2_pp.C3 = 8'd                  67;
defparam Ur3_n_2_pp.C4 = 8'd                 214;
defparam Ur3_n_2_pp.C5 = 8'd                  30;
defparam Ur3_n_2_pp.C6 = 8'd                 209;
defparam Ur3_n_2_pp.C7 = 8'd                  25;
defparam Ur3_n_2_pp.C8 = 8'd                   1;
defparam Ur3_n_2_pp.C9 = 8'd                  73;
defparam Ur3_n_2_pp.CA = 8'd                 252;
defparam Ur3_n_2_pp.CB = 8'd                  68;
defparam Ur3_n_2_pp.CC = 8'd                 215;
defparam Ur3_n_2_pp.CD = 8'd                  31;
defparam Ur3_n_2_pp.CE = 8'd                 210;
defparam Ur3_n_2_pp.CF = 8'd                  26;
assign lut_val_3_n_2_pp[13] = lut_val_3_n_2_pp[7];
assign lut_val_3_n_2_pp[12] = lut_val_3_n_2_pp[7];
assign lut_val_3_n_2_pp[11] = lut_val_3_n_2_pp[7];
assign lut_val_3_n_2_pp[10] = lut_val_3_n_2_pp[7];
assign lut_val_3_n_2_pp[9] = lut_val_3_n_2_pp[7];
assign lut_val_3_n_2_pp[8] = lut_val_3_n_2_pp[7];
wire [13:0] lut_val_3_n_3_pp;
rom_lut_r_cen Ur3_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[3],sym_res_14_n[3],sym_res_13_n[3],sym_res_12_n[3] } ), .data_out( lut_val_3_n_3_pp[7:0]) ) ;
 defparam Ur3_n_3_pp.DATA_WIDTH = 8;
defparam Ur3_n_3_pp.C0 = 8'd                   0;
defparam Ur3_n_3_pp.C1 = 8'd                  72;
defparam Ur3_n_3_pp.C2 = 8'd                 251;
defparam Ur3_n_3_pp.C3 = 8'd                  67;
defparam Ur3_n_3_pp.C4 = 8'd                 214;
defparam Ur3_n_3_pp.C5 = 8'd                  30;
defparam Ur3_n_3_pp.C6 = 8'd                 209;
defparam Ur3_n_3_pp.C7 = 8'd                  25;
defparam Ur3_n_3_pp.C8 = 8'd                   1;
defparam Ur3_n_3_pp.C9 = 8'd                  73;
defparam Ur3_n_3_pp.CA = 8'd                 252;
defparam Ur3_n_3_pp.CB = 8'd                  68;
defparam Ur3_n_3_pp.CC = 8'd                 215;
defparam Ur3_n_3_pp.CD = 8'd                  31;
defparam Ur3_n_3_pp.CE = 8'd                 210;
defparam Ur3_n_3_pp.CF = 8'd                  26;
assign lut_val_3_n_3_pp[13] = lut_val_3_n_3_pp[7];
assign lut_val_3_n_3_pp[12] = lut_val_3_n_3_pp[7];
assign lut_val_3_n_3_pp[11] = lut_val_3_n_3_pp[7];
assign lut_val_3_n_3_pp[10] = lut_val_3_n_3_pp[7];
assign lut_val_3_n_3_pp[9] = lut_val_3_n_3_pp[7];
assign lut_val_3_n_3_pp[8] = lut_val_3_n_3_pp[7];
wire [13:0] lut_val_3_n_4_pp;
rom_lut_r_cen Ur3_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[4],sym_res_14_n[4],sym_res_13_n[4],sym_res_12_n[4] } ), .data_out( lut_val_3_n_4_pp[7:0]) ) ;
 defparam Ur3_n_4_pp.DATA_WIDTH = 8;
defparam Ur3_n_4_pp.C0 = 8'd                   0;
defparam Ur3_n_4_pp.C1 = 8'd                  72;
defparam Ur3_n_4_pp.C2 = 8'd                 251;
defparam Ur3_n_4_pp.C3 = 8'd                  67;
defparam Ur3_n_4_pp.C4 = 8'd                 214;
defparam Ur3_n_4_pp.C5 = 8'd                  30;
defparam Ur3_n_4_pp.C6 = 8'd                 209;
defparam Ur3_n_4_pp.C7 = 8'd                  25;
defparam Ur3_n_4_pp.C8 = 8'd                   1;
defparam Ur3_n_4_pp.C9 = 8'd                  73;
defparam Ur3_n_4_pp.CA = 8'd                 252;
defparam Ur3_n_4_pp.CB = 8'd                  68;
defparam Ur3_n_4_pp.CC = 8'd                 215;
defparam Ur3_n_4_pp.CD = 8'd                  31;
defparam Ur3_n_4_pp.CE = 8'd                 210;
defparam Ur3_n_4_pp.CF = 8'd                  26;
assign lut_val_3_n_4_pp[13] = lut_val_3_n_4_pp[7];
assign lut_val_3_n_4_pp[12] = lut_val_3_n_4_pp[7];
assign lut_val_3_n_4_pp[11] = lut_val_3_n_4_pp[7];
assign lut_val_3_n_4_pp[10] = lut_val_3_n_4_pp[7];
assign lut_val_3_n_4_pp[9] = lut_val_3_n_4_pp[7];
assign lut_val_3_n_4_pp[8] = lut_val_3_n_4_pp[7];
wire [13:0] lut_val_3_n_5_pp;
rom_lut_r_cen Ur3_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[5],sym_res_14_n[5],sym_res_13_n[5],sym_res_12_n[5] } ), .data_out( lut_val_3_n_5_pp[7:0]) ) ;
 defparam Ur3_n_5_pp.DATA_WIDTH = 8;
defparam Ur3_n_5_pp.C0 = 8'd                   0;
defparam Ur3_n_5_pp.C1 = 8'd                  72;
defparam Ur3_n_5_pp.C2 = 8'd                 251;
defparam Ur3_n_5_pp.C3 = 8'd                  67;
defparam Ur3_n_5_pp.C4 = 8'd                 214;
defparam Ur3_n_5_pp.C5 = 8'd                  30;
defparam Ur3_n_5_pp.C6 = 8'd                 209;
defparam Ur3_n_5_pp.C7 = 8'd                  25;
defparam Ur3_n_5_pp.C8 = 8'd                   1;
defparam Ur3_n_5_pp.C9 = 8'd                  73;
defparam Ur3_n_5_pp.CA = 8'd                 252;
defparam Ur3_n_5_pp.CB = 8'd                  68;
defparam Ur3_n_5_pp.CC = 8'd                 215;
defparam Ur3_n_5_pp.CD = 8'd                  31;
defparam Ur3_n_5_pp.CE = 8'd                 210;
defparam Ur3_n_5_pp.CF = 8'd                  26;
assign lut_val_3_n_5_pp[13] = lut_val_3_n_5_pp[7];
assign lut_val_3_n_5_pp[12] = lut_val_3_n_5_pp[7];
assign lut_val_3_n_5_pp[11] = lut_val_3_n_5_pp[7];
assign lut_val_3_n_5_pp[10] = lut_val_3_n_5_pp[7];
assign lut_val_3_n_5_pp[9] = lut_val_3_n_5_pp[7];
assign lut_val_3_n_5_pp[8] = lut_val_3_n_5_pp[7];
wire [13:0] lut_val_3_n_6_pp;
rom_lut_r_cen Ur3_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[6],sym_res_14_n[6],sym_res_13_n[6],sym_res_12_n[6] } ), .data_out( lut_val_3_n_6_pp[7:0]) ) ;
 defparam Ur3_n_6_pp.DATA_WIDTH = 8;
defparam Ur3_n_6_pp.C0 = 8'd                   0;
defparam Ur3_n_6_pp.C1 = 8'd                  72;
defparam Ur3_n_6_pp.C2 = 8'd                 251;
defparam Ur3_n_6_pp.C3 = 8'd                  67;
defparam Ur3_n_6_pp.C4 = 8'd                 214;
defparam Ur3_n_6_pp.C5 = 8'd                  30;
defparam Ur3_n_6_pp.C6 = 8'd                 209;
defparam Ur3_n_6_pp.C7 = 8'd                  25;
defparam Ur3_n_6_pp.C8 = 8'd                   1;
defparam Ur3_n_6_pp.C9 = 8'd                  73;
defparam Ur3_n_6_pp.CA = 8'd                 252;
defparam Ur3_n_6_pp.CB = 8'd                  68;
defparam Ur3_n_6_pp.CC = 8'd                 215;
defparam Ur3_n_6_pp.CD = 8'd                  31;
defparam Ur3_n_6_pp.CE = 8'd                 210;
defparam Ur3_n_6_pp.CF = 8'd                  26;
assign lut_val_3_n_6_pp[13] = lut_val_3_n_6_pp[7];
assign lut_val_3_n_6_pp[12] = lut_val_3_n_6_pp[7];
assign lut_val_3_n_6_pp[11] = lut_val_3_n_6_pp[7];
assign lut_val_3_n_6_pp[10] = lut_val_3_n_6_pp[7];
assign lut_val_3_n_6_pp[9] = lut_val_3_n_6_pp[7];
assign lut_val_3_n_6_pp[8] = lut_val_3_n_6_pp[7];
wire [13:0] lut_val_3_n_7_pp;
rom_lut_r_cen Ur3_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[7],sym_res_14_n[7],sym_res_13_n[7],sym_res_12_n[7] } ), .data_out( lut_val_3_n_7_pp[7:0]) ) ;
 defparam Ur3_n_7_pp.DATA_WIDTH = 8;
defparam Ur3_n_7_pp.C0 = 8'd                   0;
defparam Ur3_n_7_pp.C1 = 8'd                  72;
defparam Ur3_n_7_pp.C2 = 8'd                 251;
defparam Ur3_n_7_pp.C3 = 8'd                  67;
defparam Ur3_n_7_pp.C4 = 8'd                 214;
defparam Ur3_n_7_pp.C5 = 8'd                  30;
defparam Ur3_n_7_pp.C6 = 8'd                 209;
defparam Ur3_n_7_pp.C7 = 8'd                  25;
defparam Ur3_n_7_pp.C8 = 8'd                   1;
defparam Ur3_n_7_pp.C9 = 8'd                  73;
defparam Ur3_n_7_pp.CA = 8'd                 252;
defparam Ur3_n_7_pp.CB = 8'd                  68;
defparam Ur3_n_7_pp.CC = 8'd                 215;
defparam Ur3_n_7_pp.CD = 8'd                  31;
defparam Ur3_n_7_pp.CE = 8'd                 210;
defparam Ur3_n_7_pp.CF = 8'd                  26;
assign lut_val_3_n_7_pp[13] = lut_val_3_n_7_pp[7];
assign lut_val_3_n_7_pp[12] = lut_val_3_n_7_pp[7];
assign lut_val_3_n_7_pp[11] = lut_val_3_n_7_pp[7];
assign lut_val_3_n_7_pp[10] = lut_val_3_n_7_pp[7];
assign lut_val_3_n_7_pp[9] = lut_val_3_n_7_pp[7];
assign lut_val_3_n_7_pp[8] = lut_val_3_n_7_pp[7];
wire [13:0] lut_val_3_n_8_pp;
rom_lut_r_cen Ur3_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[8],sym_res_14_n[8],sym_res_13_n[8],sym_res_12_n[8] } ), .data_out( lut_val_3_n_8_pp[7:0]) ) ;
 defparam Ur3_n_8_pp.DATA_WIDTH = 8;
defparam Ur3_n_8_pp.C0 = 8'd                   0;
defparam Ur3_n_8_pp.C1 = 8'd                  72;
defparam Ur3_n_8_pp.C2 = 8'd                 251;
defparam Ur3_n_8_pp.C3 = 8'd                  67;
defparam Ur3_n_8_pp.C4 = 8'd                 214;
defparam Ur3_n_8_pp.C5 = 8'd                  30;
defparam Ur3_n_8_pp.C6 = 8'd                 209;
defparam Ur3_n_8_pp.C7 = 8'd                  25;
defparam Ur3_n_8_pp.C8 = 8'd                   1;
defparam Ur3_n_8_pp.C9 = 8'd                  73;
defparam Ur3_n_8_pp.CA = 8'd                 252;
defparam Ur3_n_8_pp.CB = 8'd                  68;
defparam Ur3_n_8_pp.CC = 8'd                 215;
defparam Ur3_n_8_pp.CD = 8'd                  31;
defparam Ur3_n_8_pp.CE = 8'd                 210;
defparam Ur3_n_8_pp.CF = 8'd                  26;
assign lut_val_3_n_8_pp[13] = lut_val_3_n_8_pp[7];
assign lut_val_3_n_8_pp[12] = lut_val_3_n_8_pp[7];
assign lut_val_3_n_8_pp[11] = lut_val_3_n_8_pp[7];
assign lut_val_3_n_8_pp[10] = lut_val_3_n_8_pp[7];
assign lut_val_3_n_8_pp[9] = lut_val_3_n_8_pp[7];
assign lut_val_3_n_8_pp[8] = lut_val_3_n_8_pp[7];
wire [13:0] lut_val_3_n_9_pp;
rom_lut_r_cen Ur3_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[9],sym_res_14_n[9],sym_res_13_n[9],sym_res_12_n[9] } ), .data_out( lut_val_3_n_9_pp[7:0]) ) ;
 defparam Ur3_n_9_pp.DATA_WIDTH = 8;
defparam Ur3_n_9_pp.C0 = 8'd                   0;
defparam Ur3_n_9_pp.C1 = 8'd                  72;
defparam Ur3_n_9_pp.C2 = 8'd                 251;
defparam Ur3_n_9_pp.C3 = 8'd                  67;
defparam Ur3_n_9_pp.C4 = 8'd                 214;
defparam Ur3_n_9_pp.C5 = 8'd                  30;
defparam Ur3_n_9_pp.C6 = 8'd                 209;
defparam Ur3_n_9_pp.C7 = 8'd                  25;
defparam Ur3_n_9_pp.C8 = 8'd                   1;
defparam Ur3_n_9_pp.C9 = 8'd                  73;
defparam Ur3_n_9_pp.CA = 8'd                 252;
defparam Ur3_n_9_pp.CB = 8'd                  68;
defparam Ur3_n_9_pp.CC = 8'd                 215;
defparam Ur3_n_9_pp.CD = 8'd                  31;
defparam Ur3_n_9_pp.CE = 8'd                 210;
defparam Ur3_n_9_pp.CF = 8'd                  26;
assign lut_val_3_n_9_pp[13] = lut_val_3_n_9_pp[7];
assign lut_val_3_n_9_pp[12] = lut_val_3_n_9_pp[7];
assign lut_val_3_n_9_pp[11] = lut_val_3_n_9_pp[7];
assign lut_val_3_n_9_pp[10] = lut_val_3_n_9_pp[7];
assign lut_val_3_n_9_pp[9] = lut_val_3_n_9_pp[7];
assign lut_val_3_n_9_pp[8] = lut_val_3_n_9_pp[7];
wire [13:0] lut_val_3_n_10_pp;
rom_lut_r_cen Ur3_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[10],sym_res_14_n[10],sym_res_13_n[10],sym_res_12_n[10] } ), .data_out( lut_val_3_n_10_pp[7:0]) ) ;
 defparam Ur3_n_10_pp.DATA_WIDTH = 8;
defparam Ur3_n_10_pp.C0 = 8'd                   0;
defparam Ur3_n_10_pp.C1 = 8'd                  72;
defparam Ur3_n_10_pp.C2 = 8'd                 251;
defparam Ur3_n_10_pp.C3 = 8'd                  67;
defparam Ur3_n_10_pp.C4 = 8'd                 214;
defparam Ur3_n_10_pp.C5 = 8'd                  30;
defparam Ur3_n_10_pp.C6 = 8'd                 209;
defparam Ur3_n_10_pp.C7 = 8'd                  25;
defparam Ur3_n_10_pp.C8 = 8'd                   1;
defparam Ur3_n_10_pp.C9 = 8'd                  73;
defparam Ur3_n_10_pp.CA = 8'd                 252;
defparam Ur3_n_10_pp.CB = 8'd                  68;
defparam Ur3_n_10_pp.CC = 8'd                 215;
defparam Ur3_n_10_pp.CD = 8'd                  31;
defparam Ur3_n_10_pp.CE = 8'd                 210;
defparam Ur3_n_10_pp.CF = 8'd                  26;
assign lut_val_3_n_10_pp[13] = lut_val_3_n_10_pp[7];
assign lut_val_3_n_10_pp[12] = lut_val_3_n_10_pp[7];
assign lut_val_3_n_10_pp[11] = lut_val_3_n_10_pp[7];
assign lut_val_3_n_10_pp[10] = lut_val_3_n_10_pp[7];
assign lut_val_3_n_10_pp[9] = lut_val_3_n_10_pp[7];
assign lut_val_3_n_10_pp[8] = lut_val_3_n_10_pp[7];
wire [13:0] lut_val_3_n_11_pp;
rom_lut_r_cen Ur3_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[11],sym_res_14_n[11],sym_res_13_n[11],sym_res_12_n[11] } ), .data_out( lut_val_3_n_11_pp[7:0]) ) ;
 defparam Ur3_n_11_pp.DATA_WIDTH = 8;
defparam Ur3_n_11_pp.C0 = 8'd                   0;
defparam Ur3_n_11_pp.C1 = 8'd                  72;
defparam Ur3_n_11_pp.C2 = 8'd                 251;
defparam Ur3_n_11_pp.C3 = 8'd                  67;
defparam Ur3_n_11_pp.C4 = 8'd                 214;
defparam Ur3_n_11_pp.C5 = 8'd                  30;
defparam Ur3_n_11_pp.C6 = 8'd                 209;
defparam Ur3_n_11_pp.C7 = 8'd                  25;
defparam Ur3_n_11_pp.C8 = 8'd                   1;
defparam Ur3_n_11_pp.C9 = 8'd                  73;
defparam Ur3_n_11_pp.CA = 8'd                 252;
defparam Ur3_n_11_pp.CB = 8'd                  68;
defparam Ur3_n_11_pp.CC = 8'd                 215;
defparam Ur3_n_11_pp.CD = 8'd                  31;
defparam Ur3_n_11_pp.CE = 8'd                 210;
defparam Ur3_n_11_pp.CF = 8'd                  26;
assign lut_val_3_n_11_pp[13] = lut_val_3_n_11_pp[7];
assign lut_val_3_n_11_pp[12] = lut_val_3_n_11_pp[7];
assign lut_val_3_n_11_pp[11] = lut_val_3_n_11_pp[7];
assign lut_val_3_n_11_pp[10] = lut_val_3_n_11_pp[7];
assign lut_val_3_n_11_pp[9] = lut_val_3_n_11_pp[7];
assign lut_val_3_n_11_pp[8] = lut_val_3_n_11_pp[7];
wire [13:0] lut_val_3_n_12_pp;
rom_lut_r_cen Ur3_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[12],sym_res_14_n[12],sym_res_13_n[12],sym_res_12_n[12] } ), .data_out( lut_val_3_n_12_pp[7:0]) ) ;
 defparam Ur3_n_12_pp.DATA_WIDTH = 8;
defparam Ur3_n_12_pp.C0 = 8'd                   0;
defparam Ur3_n_12_pp.C1 = 8'd                  72;
defparam Ur3_n_12_pp.C2 = 8'd                 251;
defparam Ur3_n_12_pp.C3 = 8'd                  67;
defparam Ur3_n_12_pp.C4 = 8'd                 214;
defparam Ur3_n_12_pp.C5 = 8'd                  30;
defparam Ur3_n_12_pp.C6 = 8'd                 209;
defparam Ur3_n_12_pp.C7 = 8'd                  25;
defparam Ur3_n_12_pp.C8 = 8'd                   1;
defparam Ur3_n_12_pp.C9 = 8'd                  73;
defparam Ur3_n_12_pp.CA = 8'd                 252;
defparam Ur3_n_12_pp.CB = 8'd                  68;
defparam Ur3_n_12_pp.CC = 8'd                 215;
defparam Ur3_n_12_pp.CD = 8'd                  31;
defparam Ur3_n_12_pp.CE = 8'd                 210;
defparam Ur3_n_12_pp.CF = 8'd                  26;
assign lut_val_3_n_12_pp[13] = lut_val_3_n_12_pp[7];
assign lut_val_3_n_12_pp[12] = lut_val_3_n_12_pp[7];
assign lut_val_3_n_12_pp[11] = lut_val_3_n_12_pp[7];
assign lut_val_3_n_12_pp[10] = lut_val_3_n_12_pp[7];
assign lut_val_3_n_12_pp[9] = lut_val_3_n_12_pp[7];
assign lut_val_3_n_12_pp[8] = lut_val_3_n_12_pp[7];
wire [13:0] lut_val_3_n_13_pp;
rom_lut_r_cen Ur3_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[13],sym_res_14_n[13],sym_res_13_n[13],sym_res_12_n[13] } ), .data_out( lut_val_3_n_13_pp[7:0]) ) ;
 defparam Ur3_n_13_pp.DATA_WIDTH = 8;
defparam Ur3_n_13_pp.C0 = 8'd                   0;
defparam Ur3_n_13_pp.C1 = 8'd                  72;
defparam Ur3_n_13_pp.C2 = 8'd                 251;
defparam Ur3_n_13_pp.C3 = 8'd                  67;
defparam Ur3_n_13_pp.C4 = 8'd                 214;
defparam Ur3_n_13_pp.C5 = 8'd                  30;
defparam Ur3_n_13_pp.C6 = 8'd                 209;
defparam Ur3_n_13_pp.C7 = 8'd                  25;
defparam Ur3_n_13_pp.C8 = 8'd                   1;
defparam Ur3_n_13_pp.C9 = 8'd                  73;
defparam Ur3_n_13_pp.CA = 8'd                 252;
defparam Ur3_n_13_pp.CB = 8'd                  68;
defparam Ur3_n_13_pp.CC = 8'd                 215;
defparam Ur3_n_13_pp.CD = 8'd                  31;
defparam Ur3_n_13_pp.CE = 8'd                 210;
defparam Ur3_n_13_pp.CF = 8'd                  26;
assign lut_val_3_n_13_pp[13] = lut_val_3_n_13_pp[7];
assign lut_val_3_n_13_pp[12] = lut_val_3_n_13_pp[7];
assign lut_val_3_n_13_pp[11] = lut_val_3_n_13_pp[7];
assign lut_val_3_n_13_pp[10] = lut_val_3_n_13_pp[7];
assign lut_val_3_n_13_pp[9] = lut_val_3_n_13_pp[7];
assign lut_val_3_n_13_pp[8] = lut_val_3_n_13_pp[7];
wire [13:0] lut_val_3_n_14_pp;
rom_lut_r_cen Ur3_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[14],sym_res_14_n[14],sym_res_13_n[14],sym_res_12_n[14] } ), .data_out( lut_val_3_n_14_pp[7:0]) ) ;
 defparam Ur3_n_14_pp.DATA_WIDTH = 8;
defparam Ur3_n_14_pp.C0 = 8'd                   0;
defparam Ur3_n_14_pp.C1 = 8'd                  72;
defparam Ur3_n_14_pp.C2 = 8'd                 251;
defparam Ur3_n_14_pp.C3 = 8'd                  67;
defparam Ur3_n_14_pp.C4 = 8'd                 214;
defparam Ur3_n_14_pp.C5 = 8'd                  30;
defparam Ur3_n_14_pp.C6 = 8'd                 209;
defparam Ur3_n_14_pp.C7 = 8'd                  25;
defparam Ur3_n_14_pp.C8 = 8'd                   1;
defparam Ur3_n_14_pp.C9 = 8'd                  73;
defparam Ur3_n_14_pp.CA = 8'd                 252;
defparam Ur3_n_14_pp.CB = 8'd                  68;
defparam Ur3_n_14_pp.CC = 8'd                 215;
defparam Ur3_n_14_pp.CD = 8'd                  31;
defparam Ur3_n_14_pp.CE = 8'd                 210;
defparam Ur3_n_14_pp.CF = 8'd                  26;
assign lut_val_3_n_14_pp[13] = lut_val_3_n_14_pp[7];
assign lut_val_3_n_14_pp[12] = lut_val_3_n_14_pp[7];
assign lut_val_3_n_14_pp[11] = lut_val_3_n_14_pp[7];
assign lut_val_3_n_14_pp[10] = lut_val_3_n_14_pp[7];
assign lut_val_3_n_14_pp[9] = lut_val_3_n_14_pp[7];
assign lut_val_3_n_14_pp[8] = lut_val_3_n_14_pp[7];
wire [13:0] lut_val_3_n_15_pp;
rom_lut_r_cen Ur3_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_15_n[15],sym_res_14_n[15],sym_res_13_n[15],sym_res_12_n[15] } ), .data_out( lut_val_3_n_15_pp[7:0]) ) ;
 defparam Ur3_n_15_pp.DATA_WIDTH = 8;
defparam Ur3_n_15_pp.C0 = 8'd                   0;
defparam Ur3_n_15_pp.C1 = 8'd                  72;
defparam Ur3_n_15_pp.C2 = 8'd                 251;
defparam Ur3_n_15_pp.C3 = 8'd                  67;
defparam Ur3_n_15_pp.C4 = 8'd                 214;
defparam Ur3_n_15_pp.C5 = 8'd                  30;
defparam Ur3_n_15_pp.C6 = 8'd                 209;
defparam Ur3_n_15_pp.C7 = 8'd                  25;
defparam Ur3_n_15_pp.C8 = 8'd                   1;
defparam Ur3_n_15_pp.C9 = 8'd                  73;
defparam Ur3_n_15_pp.CA = 8'd                 252;
defparam Ur3_n_15_pp.CB = 8'd                  68;
defparam Ur3_n_15_pp.CC = 8'd                 215;
defparam Ur3_n_15_pp.CD = 8'd                  31;
defparam Ur3_n_15_pp.CE = 8'd                 210;
defparam Ur3_n_15_pp.CF = 8'd                  26;
assign lut_val_3_n_15_pp[13] = lut_val_3_n_15_pp[7];
assign lut_val_3_n_15_pp[12] = lut_val_3_n_15_pp[7];
assign lut_val_3_n_15_pp[11] = lut_val_3_n_15_pp[7];
assign lut_val_3_n_15_pp[10] = lut_val_3_n_15_pp[7];
assign lut_val_3_n_15_pp[9] = lut_val_3_n_15_pp[7];
assign lut_val_3_n_15_pp[8] = lut_val_3_n_15_pp[7];
wire [13:0] lut_val_4_n_0_pp;
rom_lut_r_cen Ur4_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[0],sym_res_18_n[0],sym_res_17_n[0],sym_res_16_n[0] } ), .data_out( lut_val_4_n_0_pp[9:0]) ) ;
 defparam Ur4_n_0_pp.DATA_WIDTH = 10;
defparam Ur4_n_0_pp.C0 = 10'd                   0;
defparam Ur4_n_0_pp.C1 = 10'd                  55;
defparam Ur4_n_0_pp.C2 = 10'd                   9;
defparam Ur4_n_0_pp.C3 = 10'd                  64;
defparam Ur4_n_0_pp.C4 = 10'd                 877;
defparam Ur4_n_0_pp.C5 = 10'd                 932;
defparam Ur4_n_0_pp.C6 = 10'd                 886;
defparam Ur4_n_0_pp.C7 = 10'd                 941;
defparam Ur4_n_0_pp.C8 = 10'd                 743;
defparam Ur4_n_0_pp.C9 = 10'd                 798;
defparam Ur4_n_0_pp.CA = 10'd                 752;
defparam Ur4_n_0_pp.CB = 10'd                 807;
defparam Ur4_n_0_pp.CC = 10'd                 596;
defparam Ur4_n_0_pp.CD = 10'd                 651;
defparam Ur4_n_0_pp.CE = 10'd                 605;
defparam Ur4_n_0_pp.CF = 10'd                 660;
assign lut_val_4_n_0_pp[13] = lut_val_4_n_0_pp[9];
assign lut_val_4_n_0_pp[12] = lut_val_4_n_0_pp[9];
assign lut_val_4_n_0_pp[11] = lut_val_4_n_0_pp[9];
assign lut_val_4_n_0_pp[10] = lut_val_4_n_0_pp[9];
wire [13:0] lut_val_4_n_1_pp;
rom_lut_r_cen Ur4_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[1],sym_res_18_n[1],sym_res_17_n[1],sym_res_16_n[1] } ), .data_out( lut_val_4_n_1_pp[9:0]) ) ;
 defparam Ur4_n_1_pp.DATA_WIDTH = 10;
defparam Ur4_n_1_pp.C0 = 10'd                   0;
defparam Ur4_n_1_pp.C1 = 10'd                  55;
defparam Ur4_n_1_pp.C2 = 10'd                   9;
defparam Ur4_n_1_pp.C3 = 10'd                  64;
defparam Ur4_n_1_pp.C4 = 10'd                 877;
defparam Ur4_n_1_pp.C5 = 10'd                 932;
defparam Ur4_n_1_pp.C6 = 10'd                 886;
defparam Ur4_n_1_pp.C7 = 10'd                 941;
defparam Ur4_n_1_pp.C8 = 10'd                 743;
defparam Ur4_n_1_pp.C9 = 10'd                 798;
defparam Ur4_n_1_pp.CA = 10'd                 752;
defparam Ur4_n_1_pp.CB = 10'd                 807;
defparam Ur4_n_1_pp.CC = 10'd                 596;
defparam Ur4_n_1_pp.CD = 10'd                 651;
defparam Ur4_n_1_pp.CE = 10'd                 605;
defparam Ur4_n_1_pp.CF = 10'd                 660;
assign lut_val_4_n_1_pp[13] = lut_val_4_n_1_pp[9];
assign lut_val_4_n_1_pp[12] = lut_val_4_n_1_pp[9];
assign lut_val_4_n_1_pp[11] = lut_val_4_n_1_pp[9];
assign lut_val_4_n_1_pp[10] = lut_val_4_n_1_pp[9];
wire [13:0] lut_val_4_n_2_pp;
rom_lut_r_cen Ur4_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[2],sym_res_18_n[2],sym_res_17_n[2],sym_res_16_n[2] } ), .data_out( lut_val_4_n_2_pp[9:0]) ) ;
 defparam Ur4_n_2_pp.DATA_WIDTH = 10;
defparam Ur4_n_2_pp.C0 = 10'd                   0;
defparam Ur4_n_2_pp.C1 = 10'd                  55;
defparam Ur4_n_2_pp.C2 = 10'd                   9;
defparam Ur4_n_2_pp.C3 = 10'd                  64;
defparam Ur4_n_2_pp.C4 = 10'd                 877;
defparam Ur4_n_2_pp.C5 = 10'd                 932;
defparam Ur4_n_2_pp.C6 = 10'd                 886;
defparam Ur4_n_2_pp.C7 = 10'd                 941;
defparam Ur4_n_2_pp.C8 = 10'd                 743;
defparam Ur4_n_2_pp.C9 = 10'd                 798;
defparam Ur4_n_2_pp.CA = 10'd                 752;
defparam Ur4_n_2_pp.CB = 10'd                 807;
defparam Ur4_n_2_pp.CC = 10'd                 596;
defparam Ur4_n_2_pp.CD = 10'd                 651;
defparam Ur4_n_2_pp.CE = 10'd                 605;
defparam Ur4_n_2_pp.CF = 10'd                 660;
assign lut_val_4_n_2_pp[13] = lut_val_4_n_2_pp[9];
assign lut_val_4_n_2_pp[12] = lut_val_4_n_2_pp[9];
assign lut_val_4_n_2_pp[11] = lut_val_4_n_2_pp[9];
assign lut_val_4_n_2_pp[10] = lut_val_4_n_2_pp[9];
wire [13:0] lut_val_4_n_3_pp;
rom_lut_r_cen Ur4_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[3],sym_res_18_n[3],sym_res_17_n[3],sym_res_16_n[3] } ), .data_out( lut_val_4_n_3_pp[9:0]) ) ;
 defparam Ur4_n_3_pp.DATA_WIDTH = 10;
defparam Ur4_n_3_pp.C0 = 10'd                   0;
defparam Ur4_n_3_pp.C1 = 10'd                  55;
defparam Ur4_n_3_pp.C2 = 10'd                   9;
defparam Ur4_n_3_pp.C3 = 10'd                  64;
defparam Ur4_n_3_pp.C4 = 10'd                 877;
defparam Ur4_n_3_pp.C5 = 10'd                 932;
defparam Ur4_n_3_pp.C6 = 10'd                 886;
defparam Ur4_n_3_pp.C7 = 10'd                 941;
defparam Ur4_n_3_pp.C8 = 10'd                 743;
defparam Ur4_n_3_pp.C9 = 10'd                 798;
defparam Ur4_n_3_pp.CA = 10'd                 752;
defparam Ur4_n_3_pp.CB = 10'd                 807;
defparam Ur4_n_3_pp.CC = 10'd                 596;
defparam Ur4_n_3_pp.CD = 10'd                 651;
defparam Ur4_n_3_pp.CE = 10'd                 605;
defparam Ur4_n_3_pp.CF = 10'd                 660;
assign lut_val_4_n_3_pp[13] = lut_val_4_n_3_pp[9];
assign lut_val_4_n_3_pp[12] = lut_val_4_n_3_pp[9];
assign lut_val_4_n_3_pp[11] = lut_val_4_n_3_pp[9];
assign lut_val_4_n_3_pp[10] = lut_val_4_n_3_pp[9];
wire [13:0] lut_val_4_n_4_pp;
rom_lut_r_cen Ur4_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[4],sym_res_18_n[4],sym_res_17_n[4],sym_res_16_n[4] } ), .data_out( lut_val_4_n_4_pp[9:0]) ) ;
 defparam Ur4_n_4_pp.DATA_WIDTH = 10;
defparam Ur4_n_4_pp.C0 = 10'd                   0;
defparam Ur4_n_4_pp.C1 = 10'd                  55;
defparam Ur4_n_4_pp.C2 = 10'd                   9;
defparam Ur4_n_4_pp.C3 = 10'd                  64;
defparam Ur4_n_4_pp.C4 = 10'd                 877;
defparam Ur4_n_4_pp.C5 = 10'd                 932;
defparam Ur4_n_4_pp.C6 = 10'd                 886;
defparam Ur4_n_4_pp.C7 = 10'd                 941;
defparam Ur4_n_4_pp.C8 = 10'd                 743;
defparam Ur4_n_4_pp.C9 = 10'd                 798;
defparam Ur4_n_4_pp.CA = 10'd                 752;
defparam Ur4_n_4_pp.CB = 10'd                 807;
defparam Ur4_n_4_pp.CC = 10'd                 596;
defparam Ur4_n_4_pp.CD = 10'd                 651;
defparam Ur4_n_4_pp.CE = 10'd                 605;
defparam Ur4_n_4_pp.CF = 10'd                 660;
assign lut_val_4_n_4_pp[13] = lut_val_4_n_4_pp[9];
assign lut_val_4_n_4_pp[12] = lut_val_4_n_4_pp[9];
assign lut_val_4_n_4_pp[11] = lut_val_4_n_4_pp[9];
assign lut_val_4_n_4_pp[10] = lut_val_4_n_4_pp[9];
wire [13:0] lut_val_4_n_5_pp;
rom_lut_r_cen Ur4_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[5],sym_res_18_n[5],sym_res_17_n[5],sym_res_16_n[5] } ), .data_out( lut_val_4_n_5_pp[9:0]) ) ;
 defparam Ur4_n_5_pp.DATA_WIDTH = 10;
defparam Ur4_n_5_pp.C0 = 10'd                   0;
defparam Ur4_n_5_pp.C1 = 10'd                  55;
defparam Ur4_n_5_pp.C2 = 10'd                   9;
defparam Ur4_n_5_pp.C3 = 10'd                  64;
defparam Ur4_n_5_pp.C4 = 10'd                 877;
defparam Ur4_n_5_pp.C5 = 10'd                 932;
defparam Ur4_n_5_pp.C6 = 10'd                 886;
defparam Ur4_n_5_pp.C7 = 10'd                 941;
defparam Ur4_n_5_pp.C8 = 10'd                 743;
defparam Ur4_n_5_pp.C9 = 10'd                 798;
defparam Ur4_n_5_pp.CA = 10'd                 752;
defparam Ur4_n_5_pp.CB = 10'd                 807;
defparam Ur4_n_5_pp.CC = 10'd                 596;
defparam Ur4_n_5_pp.CD = 10'd                 651;
defparam Ur4_n_5_pp.CE = 10'd                 605;
defparam Ur4_n_5_pp.CF = 10'd                 660;
assign lut_val_4_n_5_pp[13] = lut_val_4_n_5_pp[9];
assign lut_val_4_n_5_pp[12] = lut_val_4_n_5_pp[9];
assign lut_val_4_n_5_pp[11] = lut_val_4_n_5_pp[9];
assign lut_val_4_n_5_pp[10] = lut_val_4_n_5_pp[9];
wire [13:0] lut_val_4_n_6_pp;
rom_lut_r_cen Ur4_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[6],sym_res_18_n[6],sym_res_17_n[6],sym_res_16_n[6] } ), .data_out( lut_val_4_n_6_pp[9:0]) ) ;
 defparam Ur4_n_6_pp.DATA_WIDTH = 10;
defparam Ur4_n_6_pp.C0 = 10'd                   0;
defparam Ur4_n_6_pp.C1 = 10'd                  55;
defparam Ur4_n_6_pp.C2 = 10'd                   9;
defparam Ur4_n_6_pp.C3 = 10'd                  64;
defparam Ur4_n_6_pp.C4 = 10'd                 877;
defparam Ur4_n_6_pp.C5 = 10'd                 932;
defparam Ur4_n_6_pp.C6 = 10'd                 886;
defparam Ur4_n_6_pp.C7 = 10'd                 941;
defparam Ur4_n_6_pp.C8 = 10'd                 743;
defparam Ur4_n_6_pp.C9 = 10'd                 798;
defparam Ur4_n_6_pp.CA = 10'd                 752;
defparam Ur4_n_6_pp.CB = 10'd                 807;
defparam Ur4_n_6_pp.CC = 10'd                 596;
defparam Ur4_n_6_pp.CD = 10'd                 651;
defparam Ur4_n_6_pp.CE = 10'd                 605;
defparam Ur4_n_6_pp.CF = 10'd                 660;
assign lut_val_4_n_6_pp[13] = lut_val_4_n_6_pp[9];
assign lut_val_4_n_6_pp[12] = lut_val_4_n_6_pp[9];
assign lut_val_4_n_6_pp[11] = lut_val_4_n_6_pp[9];
assign lut_val_4_n_6_pp[10] = lut_val_4_n_6_pp[9];
wire [13:0] lut_val_4_n_7_pp;
rom_lut_r_cen Ur4_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[7],sym_res_18_n[7],sym_res_17_n[7],sym_res_16_n[7] } ), .data_out( lut_val_4_n_7_pp[9:0]) ) ;
 defparam Ur4_n_7_pp.DATA_WIDTH = 10;
defparam Ur4_n_7_pp.C0 = 10'd                   0;
defparam Ur4_n_7_pp.C1 = 10'd                  55;
defparam Ur4_n_7_pp.C2 = 10'd                   9;
defparam Ur4_n_7_pp.C3 = 10'd                  64;
defparam Ur4_n_7_pp.C4 = 10'd                 877;
defparam Ur4_n_7_pp.C5 = 10'd                 932;
defparam Ur4_n_7_pp.C6 = 10'd                 886;
defparam Ur4_n_7_pp.C7 = 10'd                 941;
defparam Ur4_n_7_pp.C8 = 10'd                 743;
defparam Ur4_n_7_pp.C9 = 10'd                 798;
defparam Ur4_n_7_pp.CA = 10'd                 752;
defparam Ur4_n_7_pp.CB = 10'd                 807;
defparam Ur4_n_7_pp.CC = 10'd                 596;
defparam Ur4_n_7_pp.CD = 10'd                 651;
defparam Ur4_n_7_pp.CE = 10'd                 605;
defparam Ur4_n_7_pp.CF = 10'd                 660;
assign lut_val_4_n_7_pp[13] = lut_val_4_n_7_pp[9];
assign lut_val_4_n_7_pp[12] = lut_val_4_n_7_pp[9];
assign lut_val_4_n_7_pp[11] = lut_val_4_n_7_pp[9];
assign lut_val_4_n_7_pp[10] = lut_val_4_n_7_pp[9];
wire [13:0] lut_val_4_n_8_pp;
rom_lut_r_cen Ur4_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[8],sym_res_18_n[8],sym_res_17_n[8],sym_res_16_n[8] } ), .data_out( lut_val_4_n_8_pp[9:0]) ) ;
 defparam Ur4_n_8_pp.DATA_WIDTH = 10;
defparam Ur4_n_8_pp.C0 = 10'd                   0;
defparam Ur4_n_8_pp.C1 = 10'd                  55;
defparam Ur4_n_8_pp.C2 = 10'd                   9;
defparam Ur4_n_8_pp.C3 = 10'd                  64;
defparam Ur4_n_8_pp.C4 = 10'd                 877;
defparam Ur4_n_8_pp.C5 = 10'd                 932;
defparam Ur4_n_8_pp.C6 = 10'd                 886;
defparam Ur4_n_8_pp.C7 = 10'd                 941;
defparam Ur4_n_8_pp.C8 = 10'd                 743;
defparam Ur4_n_8_pp.C9 = 10'd                 798;
defparam Ur4_n_8_pp.CA = 10'd                 752;
defparam Ur4_n_8_pp.CB = 10'd                 807;
defparam Ur4_n_8_pp.CC = 10'd                 596;
defparam Ur4_n_8_pp.CD = 10'd                 651;
defparam Ur4_n_8_pp.CE = 10'd                 605;
defparam Ur4_n_8_pp.CF = 10'd                 660;
assign lut_val_4_n_8_pp[13] = lut_val_4_n_8_pp[9];
assign lut_val_4_n_8_pp[12] = lut_val_4_n_8_pp[9];
assign lut_val_4_n_8_pp[11] = lut_val_4_n_8_pp[9];
assign lut_val_4_n_8_pp[10] = lut_val_4_n_8_pp[9];
wire [13:0] lut_val_4_n_9_pp;
rom_lut_r_cen Ur4_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[9],sym_res_18_n[9],sym_res_17_n[9],sym_res_16_n[9] } ), .data_out( lut_val_4_n_9_pp[9:0]) ) ;
 defparam Ur4_n_9_pp.DATA_WIDTH = 10;
defparam Ur4_n_9_pp.C0 = 10'd                   0;
defparam Ur4_n_9_pp.C1 = 10'd                  55;
defparam Ur4_n_9_pp.C2 = 10'd                   9;
defparam Ur4_n_9_pp.C3 = 10'd                  64;
defparam Ur4_n_9_pp.C4 = 10'd                 877;
defparam Ur4_n_9_pp.C5 = 10'd                 932;
defparam Ur4_n_9_pp.C6 = 10'd                 886;
defparam Ur4_n_9_pp.C7 = 10'd                 941;
defparam Ur4_n_9_pp.C8 = 10'd                 743;
defparam Ur4_n_9_pp.C9 = 10'd                 798;
defparam Ur4_n_9_pp.CA = 10'd                 752;
defparam Ur4_n_9_pp.CB = 10'd                 807;
defparam Ur4_n_9_pp.CC = 10'd                 596;
defparam Ur4_n_9_pp.CD = 10'd                 651;
defparam Ur4_n_9_pp.CE = 10'd                 605;
defparam Ur4_n_9_pp.CF = 10'd                 660;
assign lut_val_4_n_9_pp[13] = lut_val_4_n_9_pp[9];
assign lut_val_4_n_9_pp[12] = lut_val_4_n_9_pp[9];
assign lut_val_4_n_9_pp[11] = lut_val_4_n_9_pp[9];
assign lut_val_4_n_9_pp[10] = lut_val_4_n_9_pp[9];
wire [13:0] lut_val_4_n_10_pp;
rom_lut_r_cen Ur4_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[10],sym_res_18_n[10],sym_res_17_n[10],sym_res_16_n[10] } ), .data_out( lut_val_4_n_10_pp[9:0]) ) ;
 defparam Ur4_n_10_pp.DATA_WIDTH = 10;
defparam Ur4_n_10_pp.C0 = 10'd                   0;
defparam Ur4_n_10_pp.C1 = 10'd                  55;
defparam Ur4_n_10_pp.C2 = 10'd                   9;
defparam Ur4_n_10_pp.C3 = 10'd                  64;
defparam Ur4_n_10_pp.C4 = 10'd                 877;
defparam Ur4_n_10_pp.C5 = 10'd                 932;
defparam Ur4_n_10_pp.C6 = 10'd                 886;
defparam Ur4_n_10_pp.C7 = 10'd                 941;
defparam Ur4_n_10_pp.C8 = 10'd                 743;
defparam Ur4_n_10_pp.C9 = 10'd                 798;
defparam Ur4_n_10_pp.CA = 10'd                 752;
defparam Ur4_n_10_pp.CB = 10'd                 807;
defparam Ur4_n_10_pp.CC = 10'd                 596;
defparam Ur4_n_10_pp.CD = 10'd                 651;
defparam Ur4_n_10_pp.CE = 10'd                 605;
defparam Ur4_n_10_pp.CF = 10'd                 660;
assign lut_val_4_n_10_pp[13] = lut_val_4_n_10_pp[9];
assign lut_val_4_n_10_pp[12] = lut_val_4_n_10_pp[9];
assign lut_val_4_n_10_pp[11] = lut_val_4_n_10_pp[9];
assign lut_val_4_n_10_pp[10] = lut_val_4_n_10_pp[9];
wire [13:0] lut_val_4_n_11_pp;
rom_lut_r_cen Ur4_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[11],sym_res_18_n[11],sym_res_17_n[11],sym_res_16_n[11] } ), .data_out( lut_val_4_n_11_pp[9:0]) ) ;
 defparam Ur4_n_11_pp.DATA_WIDTH = 10;
defparam Ur4_n_11_pp.C0 = 10'd                   0;
defparam Ur4_n_11_pp.C1 = 10'd                  55;
defparam Ur4_n_11_pp.C2 = 10'd                   9;
defparam Ur4_n_11_pp.C3 = 10'd                  64;
defparam Ur4_n_11_pp.C4 = 10'd                 877;
defparam Ur4_n_11_pp.C5 = 10'd                 932;
defparam Ur4_n_11_pp.C6 = 10'd                 886;
defparam Ur4_n_11_pp.C7 = 10'd                 941;
defparam Ur4_n_11_pp.C8 = 10'd                 743;
defparam Ur4_n_11_pp.C9 = 10'd                 798;
defparam Ur4_n_11_pp.CA = 10'd                 752;
defparam Ur4_n_11_pp.CB = 10'd                 807;
defparam Ur4_n_11_pp.CC = 10'd                 596;
defparam Ur4_n_11_pp.CD = 10'd                 651;
defparam Ur4_n_11_pp.CE = 10'd                 605;
defparam Ur4_n_11_pp.CF = 10'd                 660;
assign lut_val_4_n_11_pp[13] = lut_val_4_n_11_pp[9];
assign lut_val_4_n_11_pp[12] = lut_val_4_n_11_pp[9];
assign lut_val_4_n_11_pp[11] = lut_val_4_n_11_pp[9];
assign lut_val_4_n_11_pp[10] = lut_val_4_n_11_pp[9];
wire [13:0] lut_val_4_n_12_pp;
rom_lut_r_cen Ur4_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[12],sym_res_18_n[12],sym_res_17_n[12],sym_res_16_n[12] } ), .data_out( lut_val_4_n_12_pp[9:0]) ) ;
 defparam Ur4_n_12_pp.DATA_WIDTH = 10;
defparam Ur4_n_12_pp.C0 = 10'd                   0;
defparam Ur4_n_12_pp.C1 = 10'd                  55;
defparam Ur4_n_12_pp.C2 = 10'd                   9;
defparam Ur4_n_12_pp.C3 = 10'd                  64;
defparam Ur4_n_12_pp.C4 = 10'd                 877;
defparam Ur4_n_12_pp.C5 = 10'd                 932;
defparam Ur4_n_12_pp.C6 = 10'd                 886;
defparam Ur4_n_12_pp.C7 = 10'd                 941;
defparam Ur4_n_12_pp.C8 = 10'd                 743;
defparam Ur4_n_12_pp.C9 = 10'd                 798;
defparam Ur4_n_12_pp.CA = 10'd                 752;
defparam Ur4_n_12_pp.CB = 10'd                 807;
defparam Ur4_n_12_pp.CC = 10'd                 596;
defparam Ur4_n_12_pp.CD = 10'd                 651;
defparam Ur4_n_12_pp.CE = 10'd                 605;
defparam Ur4_n_12_pp.CF = 10'd                 660;
assign lut_val_4_n_12_pp[13] = lut_val_4_n_12_pp[9];
assign lut_val_4_n_12_pp[12] = lut_val_4_n_12_pp[9];
assign lut_val_4_n_12_pp[11] = lut_val_4_n_12_pp[9];
assign lut_val_4_n_12_pp[10] = lut_val_4_n_12_pp[9];
wire [13:0] lut_val_4_n_13_pp;
rom_lut_r_cen Ur4_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[13],sym_res_18_n[13],sym_res_17_n[13],sym_res_16_n[13] } ), .data_out( lut_val_4_n_13_pp[9:0]) ) ;
 defparam Ur4_n_13_pp.DATA_WIDTH = 10;
defparam Ur4_n_13_pp.C0 = 10'd                   0;
defparam Ur4_n_13_pp.C1 = 10'd                  55;
defparam Ur4_n_13_pp.C2 = 10'd                   9;
defparam Ur4_n_13_pp.C3 = 10'd                  64;
defparam Ur4_n_13_pp.C4 = 10'd                 877;
defparam Ur4_n_13_pp.C5 = 10'd                 932;
defparam Ur4_n_13_pp.C6 = 10'd                 886;
defparam Ur4_n_13_pp.C7 = 10'd                 941;
defparam Ur4_n_13_pp.C8 = 10'd                 743;
defparam Ur4_n_13_pp.C9 = 10'd                 798;
defparam Ur4_n_13_pp.CA = 10'd                 752;
defparam Ur4_n_13_pp.CB = 10'd                 807;
defparam Ur4_n_13_pp.CC = 10'd                 596;
defparam Ur4_n_13_pp.CD = 10'd                 651;
defparam Ur4_n_13_pp.CE = 10'd                 605;
defparam Ur4_n_13_pp.CF = 10'd                 660;
assign lut_val_4_n_13_pp[13] = lut_val_4_n_13_pp[9];
assign lut_val_4_n_13_pp[12] = lut_val_4_n_13_pp[9];
assign lut_val_4_n_13_pp[11] = lut_val_4_n_13_pp[9];
assign lut_val_4_n_13_pp[10] = lut_val_4_n_13_pp[9];
wire [13:0] lut_val_4_n_14_pp;
rom_lut_r_cen Ur4_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[14],sym_res_18_n[14],sym_res_17_n[14],sym_res_16_n[14] } ), .data_out( lut_val_4_n_14_pp[9:0]) ) ;
 defparam Ur4_n_14_pp.DATA_WIDTH = 10;
defparam Ur4_n_14_pp.C0 = 10'd                   0;
defparam Ur4_n_14_pp.C1 = 10'd                  55;
defparam Ur4_n_14_pp.C2 = 10'd                   9;
defparam Ur4_n_14_pp.C3 = 10'd                  64;
defparam Ur4_n_14_pp.C4 = 10'd                 877;
defparam Ur4_n_14_pp.C5 = 10'd                 932;
defparam Ur4_n_14_pp.C6 = 10'd                 886;
defparam Ur4_n_14_pp.C7 = 10'd                 941;
defparam Ur4_n_14_pp.C8 = 10'd                 743;
defparam Ur4_n_14_pp.C9 = 10'd                 798;
defparam Ur4_n_14_pp.CA = 10'd                 752;
defparam Ur4_n_14_pp.CB = 10'd                 807;
defparam Ur4_n_14_pp.CC = 10'd                 596;
defparam Ur4_n_14_pp.CD = 10'd                 651;
defparam Ur4_n_14_pp.CE = 10'd                 605;
defparam Ur4_n_14_pp.CF = 10'd                 660;
assign lut_val_4_n_14_pp[13] = lut_val_4_n_14_pp[9];
assign lut_val_4_n_14_pp[12] = lut_val_4_n_14_pp[9];
assign lut_val_4_n_14_pp[11] = lut_val_4_n_14_pp[9];
assign lut_val_4_n_14_pp[10] = lut_val_4_n_14_pp[9];
wire [13:0] lut_val_4_n_15_pp;
rom_lut_r_cen Ur4_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_19_n[15],sym_res_18_n[15],sym_res_17_n[15],sym_res_16_n[15] } ), .data_out( lut_val_4_n_15_pp[9:0]) ) ;
 defparam Ur4_n_15_pp.DATA_WIDTH = 10;
defparam Ur4_n_15_pp.C0 = 10'd                   0;
defparam Ur4_n_15_pp.C1 = 10'd                  55;
defparam Ur4_n_15_pp.C2 = 10'd                   9;
defparam Ur4_n_15_pp.C3 = 10'd                  64;
defparam Ur4_n_15_pp.C4 = 10'd                 877;
defparam Ur4_n_15_pp.C5 = 10'd                 932;
defparam Ur4_n_15_pp.C6 = 10'd                 886;
defparam Ur4_n_15_pp.C7 = 10'd                 941;
defparam Ur4_n_15_pp.C8 = 10'd                 743;
defparam Ur4_n_15_pp.C9 = 10'd                 798;
defparam Ur4_n_15_pp.CA = 10'd                 752;
defparam Ur4_n_15_pp.CB = 10'd                 807;
defparam Ur4_n_15_pp.CC = 10'd                 596;
defparam Ur4_n_15_pp.CD = 10'd                 651;
defparam Ur4_n_15_pp.CE = 10'd                 605;
defparam Ur4_n_15_pp.CF = 10'd                 660;
assign lut_val_4_n_15_pp[13] = lut_val_4_n_15_pp[9];
assign lut_val_4_n_15_pp[12] = lut_val_4_n_15_pp[9];
assign lut_val_4_n_15_pp[11] = lut_val_4_n_15_pp[9];
assign lut_val_4_n_15_pp[10] = lut_val_4_n_15_pp[9];
wire [13:0] lut_val_5_n_0_pp;
rom_lut_r_cen Ur5_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[0],sym_res_22_n[0],sym_res_21_n[0],sym_res_20_n[0] } ), .data_out( lut_val_5_n_0_pp[9:0]) ) ;
 defparam Ur5_n_0_pp.DATA_WIDTH = 10;
defparam Ur5_n_0_pp.C0 = 10'd                   0;
defparam Ur5_n_0_pp.C1 = 10'd                 782;
defparam Ur5_n_0_pp.C2 = 10'd                 974;
defparam Ur5_n_0_pp.C3 = 10'd                 732;
defparam Ur5_n_0_pp.C4 = 10'd                 100;
defparam Ur5_n_0_pp.C5 = 10'd                 882;
defparam Ur5_n_0_pp.C6 = 10'd                  50;
defparam Ur5_n_0_pp.C7 = 10'd                 832;
defparam Ur5_n_0_pp.C8 = 10'd                  51;
defparam Ur5_n_0_pp.C9 = 10'd                 833;
defparam Ur5_n_0_pp.CA = 10'd                   1;
defparam Ur5_n_0_pp.CB = 10'd                 783;
defparam Ur5_n_0_pp.CC = 10'd                 151;
defparam Ur5_n_0_pp.CD = 10'd                 933;
defparam Ur5_n_0_pp.CE = 10'd                 101;
defparam Ur5_n_0_pp.CF = 10'd                 883;
assign lut_val_5_n_0_pp[13] = lut_val_5_n_0_pp[9];
assign lut_val_5_n_0_pp[12] = lut_val_5_n_0_pp[9];
assign lut_val_5_n_0_pp[11] = lut_val_5_n_0_pp[9];
assign lut_val_5_n_0_pp[10] = lut_val_5_n_0_pp[9];
wire [13:0] lut_val_5_n_1_pp;
rom_lut_r_cen Ur5_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[1],sym_res_22_n[1],sym_res_21_n[1],sym_res_20_n[1] } ), .data_out( lut_val_5_n_1_pp[9:0]) ) ;
 defparam Ur5_n_1_pp.DATA_WIDTH = 10;
defparam Ur5_n_1_pp.C0 = 10'd                   0;
defparam Ur5_n_1_pp.C1 = 10'd                 782;
defparam Ur5_n_1_pp.C2 = 10'd                 974;
defparam Ur5_n_1_pp.C3 = 10'd                 732;
defparam Ur5_n_1_pp.C4 = 10'd                 100;
defparam Ur5_n_1_pp.C5 = 10'd                 882;
defparam Ur5_n_1_pp.C6 = 10'd                  50;
defparam Ur5_n_1_pp.C7 = 10'd                 832;
defparam Ur5_n_1_pp.C8 = 10'd                  51;
defparam Ur5_n_1_pp.C9 = 10'd                 833;
defparam Ur5_n_1_pp.CA = 10'd                   1;
defparam Ur5_n_1_pp.CB = 10'd                 783;
defparam Ur5_n_1_pp.CC = 10'd                 151;
defparam Ur5_n_1_pp.CD = 10'd                 933;
defparam Ur5_n_1_pp.CE = 10'd                 101;
defparam Ur5_n_1_pp.CF = 10'd                 883;
assign lut_val_5_n_1_pp[13] = lut_val_5_n_1_pp[9];
assign lut_val_5_n_1_pp[12] = lut_val_5_n_1_pp[9];
assign lut_val_5_n_1_pp[11] = lut_val_5_n_1_pp[9];
assign lut_val_5_n_1_pp[10] = lut_val_5_n_1_pp[9];
wire [13:0] lut_val_5_n_2_pp;
rom_lut_r_cen Ur5_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[2],sym_res_22_n[2],sym_res_21_n[2],sym_res_20_n[2] } ), .data_out( lut_val_5_n_2_pp[9:0]) ) ;
 defparam Ur5_n_2_pp.DATA_WIDTH = 10;
defparam Ur5_n_2_pp.C0 = 10'd                   0;
defparam Ur5_n_2_pp.C1 = 10'd                 782;
defparam Ur5_n_2_pp.C2 = 10'd                 974;
defparam Ur5_n_2_pp.C3 = 10'd                 732;
defparam Ur5_n_2_pp.C4 = 10'd                 100;
defparam Ur5_n_2_pp.C5 = 10'd                 882;
defparam Ur5_n_2_pp.C6 = 10'd                  50;
defparam Ur5_n_2_pp.C7 = 10'd                 832;
defparam Ur5_n_2_pp.C8 = 10'd                  51;
defparam Ur5_n_2_pp.C9 = 10'd                 833;
defparam Ur5_n_2_pp.CA = 10'd                   1;
defparam Ur5_n_2_pp.CB = 10'd                 783;
defparam Ur5_n_2_pp.CC = 10'd                 151;
defparam Ur5_n_2_pp.CD = 10'd                 933;
defparam Ur5_n_2_pp.CE = 10'd                 101;
defparam Ur5_n_2_pp.CF = 10'd                 883;
assign lut_val_5_n_2_pp[13] = lut_val_5_n_2_pp[9];
assign lut_val_5_n_2_pp[12] = lut_val_5_n_2_pp[9];
assign lut_val_5_n_2_pp[11] = lut_val_5_n_2_pp[9];
assign lut_val_5_n_2_pp[10] = lut_val_5_n_2_pp[9];
wire [13:0] lut_val_5_n_3_pp;
rom_lut_r_cen Ur5_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[3],sym_res_22_n[3],sym_res_21_n[3],sym_res_20_n[3] } ), .data_out( lut_val_5_n_3_pp[9:0]) ) ;
 defparam Ur5_n_3_pp.DATA_WIDTH = 10;
defparam Ur5_n_3_pp.C0 = 10'd                   0;
defparam Ur5_n_3_pp.C1 = 10'd                 782;
defparam Ur5_n_3_pp.C2 = 10'd                 974;
defparam Ur5_n_3_pp.C3 = 10'd                 732;
defparam Ur5_n_3_pp.C4 = 10'd                 100;
defparam Ur5_n_3_pp.C5 = 10'd                 882;
defparam Ur5_n_3_pp.C6 = 10'd                  50;
defparam Ur5_n_3_pp.C7 = 10'd                 832;
defparam Ur5_n_3_pp.C8 = 10'd                  51;
defparam Ur5_n_3_pp.C9 = 10'd                 833;
defparam Ur5_n_3_pp.CA = 10'd                   1;
defparam Ur5_n_3_pp.CB = 10'd                 783;
defparam Ur5_n_3_pp.CC = 10'd                 151;
defparam Ur5_n_3_pp.CD = 10'd                 933;
defparam Ur5_n_3_pp.CE = 10'd                 101;
defparam Ur5_n_3_pp.CF = 10'd                 883;
assign lut_val_5_n_3_pp[13] = lut_val_5_n_3_pp[9];
assign lut_val_5_n_3_pp[12] = lut_val_5_n_3_pp[9];
assign lut_val_5_n_3_pp[11] = lut_val_5_n_3_pp[9];
assign lut_val_5_n_3_pp[10] = lut_val_5_n_3_pp[9];
wire [13:0] lut_val_5_n_4_pp;
rom_lut_r_cen Ur5_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[4],sym_res_22_n[4],sym_res_21_n[4],sym_res_20_n[4] } ), .data_out( lut_val_5_n_4_pp[9:0]) ) ;
 defparam Ur5_n_4_pp.DATA_WIDTH = 10;
defparam Ur5_n_4_pp.C0 = 10'd                   0;
defparam Ur5_n_4_pp.C1 = 10'd                 782;
defparam Ur5_n_4_pp.C2 = 10'd                 974;
defparam Ur5_n_4_pp.C3 = 10'd                 732;
defparam Ur5_n_4_pp.C4 = 10'd                 100;
defparam Ur5_n_4_pp.C5 = 10'd                 882;
defparam Ur5_n_4_pp.C6 = 10'd                  50;
defparam Ur5_n_4_pp.C7 = 10'd                 832;
defparam Ur5_n_4_pp.C8 = 10'd                  51;
defparam Ur5_n_4_pp.C9 = 10'd                 833;
defparam Ur5_n_4_pp.CA = 10'd                   1;
defparam Ur5_n_4_pp.CB = 10'd                 783;
defparam Ur5_n_4_pp.CC = 10'd                 151;
defparam Ur5_n_4_pp.CD = 10'd                 933;
defparam Ur5_n_4_pp.CE = 10'd                 101;
defparam Ur5_n_4_pp.CF = 10'd                 883;
assign lut_val_5_n_4_pp[13] = lut_val_5_n_4_pp[9];
assign lut_val_5_n_4_pp[12] = lut_val_5_n_4_pp[9];
assign lut_val_5_n_4_pp[11] = lut_val_5_n_4_pp[9];
assign lut_val_5_n_4_pp[10] = lut_val_5_n_4_pp[9];
wire [13:0] lut_val_5_n_5_pp;
rom_lut_r_cen Ur5_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[5],sym_res_22_n[5],sym_res_21_n[5],sym_res_20_n[5] } ), .data_out( lut_val_5_n_5_pp[9:0]) ) ;
 defparam Ur5_n_5_pp.DATA_WIDTH = 10;
defparam Ur5_n_5_pp.C0 = 10'd                   0;
defparam Ur5_n_5_pp.C1 = 10'd                 782;
defparam Ur5_n_5_pp.C2 = 10'd                 974;
defparam Ur5_n_5_pp.C3 = 10'd                 732;
defparam Ur5_n_5_pp.C4 = 10'd                 100;
defparam Ur5_n_5_pp.C5 = 10'd                 882;
defparam Ur5_n_5_pp.C6 = 10'd                  50;
defparam Ur5_n_5_pp.C7 = 10'd                 832;
defparam Ur5_n_5_pp.C8 = 10'd                  51;
defparam Ur5_n_5_pp.C9 = 10'd                 833;
defparam Ur5_n_5_pp.CA = 10'd                   1;
defparam Ur5_n_5_pp.CB = 10'd                 783;
defparam Ur5_n_5_pp.CC = 10'd                 151;
defparam Ur5_n_5_pp.CD = 10'd                 933;
defparam Ur5_n_5_pp.CE = 10'd                 101;
defparam Ur5_n_5_pp.CF = 10'd                 883;
assign lut_val_5_n_5_pp[13] = lut_val_5_n_5_pp[9];
assign lut_val_5_n_5_pp[12] = lut_val_5_n_5_pp[9];
assign lut_val_5_n_5_pp[11] = lut_val_5_n_5_pp[9];
assign lut_val_5_n_5_pp[10] = lut_val_5_n_5_pp[9];
wire [13:0] lut_val_5_n_6_pp;
rom_lut_r_cen Ur5_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[6],sym_res_22_n[6],sym_res_21_n[6],sym_res_20_n[6] } ), .data_out( lut_val_5_n_6_pp[9:0]) ) ;
 defparam Ur5_n_6_pp.DATA_WIDTH = 10;
defparam Ur5_n_6_pp.C0 = 10'd                   0;
defparam Ur5_n_6_pp.C1 = 10'd                 782;
defparam Ur5_n_6_pp.C2 = 10'd                 974;
defparam Ur5_n_6_pp.C3 = 10'd                 732;
defparam Ur5_n_6_pp.C4 = 10'd                 100;
defparam Ur5_n_6_pp.C5 = 10'd                 882;
defparam Ur5_n_6_pp.C6 = 10'd                  50;
defparam Ur5_n_6_pp.C7 = 10'd                 832;
defparam Ur5_n_6_pp.C8 = 10'd                  51;
defparam Ur5_n_6_pp.C9 = 10'd                 833;
defparam Ur5_n_6_pp.CA = 10'd                   1;
defparam Ur5_n_6_pp.CB = 10'd                 783;
defparam Ur5_n_6_pp.CC = 10'd                 151;
defparam Ur5_n_6_pp.CD = 10'd                 933;
defparam Ur5_n_6_pp.CE = 10'd                 101;
defparam Ur5_n_6_pp.CF = 10'd                 883;
assign lut_val_5_n_6_pp[13] = lut_val_5_n_6_pp[9];
assign lut_val_5_n_6_pp[12] = lut_val_5_n_6_pp[9];
assign lut_val_5_n_6_pp[11] = lut_val_5_n_6_pp[9];
assign lut_val_5_n_6_pp[10] = lut_val_5_n_6_pp[9];
wire [13:0] lut_val_5_n_7_pp;
rom_lut_r_cen Ur5_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[7],sym_res_22_n[7],sym_res_21_n[7],sym_res_20_n[7] } ), .data_out( lut_val_5_n_7_pp[9:0]) ) ;
 defparam Ur5_n_7_pp.DATA_WIDTH = 10;
defparam Ur5_n_7_pp.C0 = 10'd                   0;
defparam Ur5_n_7_pp.C1 = 10'd                 782;
defparam Ur5_n_7_pp.C2 = 10'd                 974;
defparam Ur5_n_7_pp.C3 = 10'd                 732;
defparam Ur5_n_7_pp.C4 = 10'd                 100;
defparam Ur5_n_7_pp.C5 = 10'd                 882;
defparam Ur5_n_7_pp.C6 = 10'd                  50;
defparam Ur5_n_7_pp.C7 = 10'd                 832;
defparam Ur5_n_7_pp.C8 = 10'd                  51;
defparam Ur5_n_7_pp.C9 = 10'd                 833;
defparam Ur5_n_7_pp.CA = 10'd                   1;
defparam Ur5_n_7_pp.CB = 10'd                 783;
defparam Ur5_n_7_pp.CC = 10'd                 151;
defparam Ur5_n_7_pp.CD = 10'd                 933;
defparam Ur5_n_7_pp.CE = 10'd                 101;
defparam Ur5_n_7_pp.CF = 10'd                 883;
assign lut_val_5_n_7_pp[13] = lut_val_5_n_7_pp[9];
assign lut_val_5_n_7_pp[12] = lut_val_5_n_7_pp[9];
assign lut_val_5_n_7_pp[11] = lut_val_5_n_7_pp[9];
assign lut_val_5_n_7_pp[10] = lut_val_5_n_7_pp[9];
wire [13:0] lut_val_5_n_8_pp;
rom_lut_r_cen Ur5_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[8],sym_res_22_n[8],sym_res_21_n[8],sym_res_20_n[8] } ), .data_out( lut_val_5_n_8_pp[9:0]) ) ;
 defparam Ur5_n_8_pp.DATA_WIDTH = 10;
defparam Ur5_n_8_pp.C0 = 10'd                   0;
defparam Ur5_n_8_pp.C1 = 10'd                 782;
defparam Ur5_n_8_pp.C2 = 10'd                 974;
defparam Ur5_n_8_pp.C3 = 10'd                 732;
defparam Ur5_n_8_pp.C4 = 10'd                 100;
defparam Ur5_n_8_pp.C5 = 10'd                 882;
defparam Ur5_n_8_pp.C6 = 10'd                  50;
defparam Ur5_n_8_pp.C7 = 10'd                 832;
defparam Ur5_n_8_pp.C8 = 10'd                  51;
defparam Ur5_n_8_pp.C9 = 10'd                 833;
defparam Ur5_n_8_pp.CA = 10'd                   1;
defparam Ur5_n_8_pp.CB = 10'd                 783;
defparam Ur5_n_8_pp.CC = 10'd                 151;
defparam Ur5_n_8_pp.CD = 10'd                 933;
defparam Ur5_n_8_pp.CE = 10'd                 101;
defparam Ur5_n_8_pp.CF = 10'd                 883;
assign lut_val_5_n_8_pp[13] = lut_val_5_n_8_pp[9];
assign lut_val_5_n_8_pp[12] = lut_val_5_n_8_pp[9];
assign lut_val_5_n_8_pp[11] = lut_val_5_n_8_pp[9];
assign lut_val_5_n_8_pp[10] = lut_val_5_n_8_pp[9];
wire [13:0] lut_val_5_n_9_pp;
rom_lut_r_cen Ur5_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[9],sym_res_22_n[9],sym_res_21_n[9],sym_res_20_n[9] } ), .data_out( lut_val_5_n_9_pp[9:0]) ) ;
 defparam Ur5_n_9_pp.DATA_WIDTH = 10;
defparam Ur5_n_9_pp.C0 = 10'd                   0;
defparam Ur5_n_9_pp.C1 = 10'd                 782;
defparam Ur5_n_9_pp.C2 = 10'd                 974;
defparam Ur5_n_9_pp.C3 = 10'd                 732;
defparam Ur5_n_9_pp.C4 = 10'd                 100;
defparam Ur5_n_9_pp.C5 = 10'd                 882;
defparam Ur5_n_9_pp.C6 = 10'd                  50;
defparam Ur5_n_9_pp.C7 = 10'd                 832;
defparam Ur5_n_9_pp.C8 = 10'd                  51;
defparam Ur5_n_9_pp.C9 = 10'd                 833;
defparam Ur5_n_9_pp.CA = 10'd                   1;
defparam Ur5_n_9_pp.CB = 10'd                 783;
defparam Ur5_n_9_pp.CC = 10'd                 151;
defparam Ur5_n_9_pp.CD = 10'd                 933;
defparam Ur5_n_9_pp.CE = 10'd                 101;
defparam Ur5_n_9_pp.CF = 10'd                 883;
assign lut_val_5_n_9_pp[13] = lut_val_5_n_9_pp[9];
assign lut_val_5_n_9_pp[12] = lut_val_5_n_9_pp[9];
assign lut_val_5_n_9_pp[11] = lut_val_5_n_9_pp[9];
assign lut_val_5_n_9_pp[10] = lut_val_5_n_9_pp[9];
wire [13:0] lut_val_5_n_10_pp;
rom_lut_r_cen Ur5_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[10],sym_res_22_n[10],sym_res_21_n[10],sym_res_20_n[10] } ), .data_out( lut_val_5_n_10_pp[9:0]) ) ;
 defparam Ur5_n_10_pp.DATA_WIDTH = 10;
defparam Ur5_n_10_pp.C0 = 10'd                   0;
defparam Ur5_n_10_pp.C1 = 10'd                 782;
defparam Ur5_n_10_pp.C2 = 10'd                 974;
defparam Ur5_n_10_pp.C3 = 10'd                 732;
defparam Ur5_n_10_pp.C4 = 10'd                 100;
defparam Ur5_n_10_pp.C5 = 10'd                 882;
defparam Ur5_n_10_pp.C6 = 10'd                  50;
defparam Ur5_n_10_pp.C7 = 10'd                 832;
defparam Ur5_n_10_pp.C8 = 10'd                  51;
defparam Ur5_n_10_pp.C9 = 10'd                 833;
defparam Ur5_n_10_pp.CA = 10'd                   1;
defparam Ur5_n_10_pp.CB = 10'd                 783;
defparam Ur5_n_10_pp.CC = 10'd                 151;
defparam Ur5_n_10_pp.CD = 10'd                 933;
defparam Ur5_n_10_pp.CE = 10'd                 101;
defparam Ur5_n_10_pp.CF = 10'd                 883;
assign lut_val_5_n_10_pp[13] = lut_val_5_n_10_pp[9];
assign lut_val_5_n_10_pp[12] = lut_val_5_n_10_pp[9];
assign lut_val_5_n_10_pp[11] = lut_val_5_n_10_pp[9];
assign lut_val_5_n_10_pp[10] = lut_val_5_n_10_pp[9];
wire [13:0] lut_val_5_n_11_pp;
rom_lut_r_cen Ur5_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[11],sym_res_22_n[11],sym_res_21_n[11],sym_res_20_n[11] } ), .data_out( lut_val_5_n_11_pp[9:0]) ) ;
 defparam Ur5_n_11_pp.DATA_WIDTH = 10;
defparam Ur5_n_11_pp.C0 = 10'd                   0;
defparam Ur5_n_11_pp.C1 = 10'd                 782;
defparam Ur5_n_11_pp.C2 = 10'd                 974;
defparam Ur5_n_11_pp.C3 = 10'd                 732;
defparam Ur5_n_11_pp.C4 = 10'd                 100;
defparam Ur5_n_11_pp.C5 = 10'd                 882;
defparam Ur5_n_11_pp.C6 = 10'd                  50;
defparam Ur5_n_11_pp.C7 = 10'd                 832;
defparam Ur5_n_11_pp.C8 = 10'd                  51;
defparam Ur5_n_11_pp.C9 = 10'd                 833;
defparam Ur5_n_11_pp.CA = 10'd                   1;
defparam Ur5_n_11_pp.CB = 10'd                 783;
defparam Ur5_n_11_pp.CC = 10'd                 151;
defparam Ur5_n_11_pp.CD = 10'd                 933;
defparam Ur5_n_11_pp.CE = 10'd                 101;
defparam Ur5_n_11_pp.CF = 10'd                 883;
assign lut_val_5_n_11_pp[13] = lut_val_5_n_11_pp[9];
assign lut_val_5_n_11_pp[12] = lut_val_5_n_11_pp[9];
assign lut_val_5_n_11_pp[11] = lut_val_5_n_11_pp[9];
assign lut_val_5_n_11_pp[10] = lut_val_5_n_11_pp[9];
wire [13:0] lut_val_5_n_12_pp;
rom_lut_r_cen Ur5_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[12],sym_res_22_n[12],sym_res_21_n[12],sym_res_20_n[12] } ), .data_out( lut_val_5_n_12_pp[9:0]) ) ;
 defparam Ur5_n_12_pp.DATA_WIDTH = 10;
defparam Ur5_n_12_pp.C0 = 10'd                   0;
defparam Ur5_n_12_pp.C1 = 10'd                 782;
defparam Ur5_n_12_pp.C2 = 10'd                 974;
defparam Ur5_n_12_pp.C3 = 10'd                 732;
defparam Ur5_n_12_pp.C4 = 10'd                 100;
defparam Ur5_n_12_pp.C5 = 10'd                 882;
defparam Ur5_n_12_pp.C6 = 10'd                  50;
defparam Ur5_n_12_pp.C7 = 10'd                 832;
defparam Ur5_n_12_pp.C8 = 10'd                  51;
defparam Ur5_n_12_pp.C9 = 10'd                 833;
defparam Ur5_n_12_pp.CA = 10'd                   1;
defparam Ur5_n_12_pp.CB = 10'd                 783;
defparam Ur5_n_12_pp.CC = 10'd                 151;
defparam Ur5_n_12_pp.CD = 10'd                 933;
defparam Ur5_n_12_pp.CE = 10'd                 101;
defparam Ur5_n_12_pp.CF = 10'd                 883;
assign lut_val_5_n_12_pp[13] = lut_val_5_n_12_pp[9];
assign lut_val_5_n_12_pp[12] = lut_val_5_n_12_pp[9];
assign lut_val_5_n_12_pp[11] = lut_val_5_n_12_pp[9];
assign lut_val_5_n_12_pp[10] = lut_val_5_n_12_pp[9];
wire [13:0] lut_val_5_n_13_pp;
rom_lut_r_cen Ur5_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[13],sym_res_22_n[13],sym_res_21_n[13],sym_res_20_n[13] } ), .data_out( lut_val_5_n_13_pp[9:0]) ) ;
 defparam Ur5_n_13_pp.DATA_WIDTH = 10;
defparam Ur5_n_13_pp.C0 = 10'd                   0;
defparam Ur5_n_13_pp.C1 = 10'd                 782;
defparam Ur5_n_13_pp.C2 = 10'd                 974;
defparam Ur5_n_13_pp.C3 = 10'd                 732;
defparam Ur5_n_13_pp.C4 = 10'd                 100;
defparam Ur5_n_13_pp.C5 = 10'd                 882;
defparam Ur5_n_13_pp.C6 = 10'd                  50;
defparam Ur5_n_13_pp.C7 = 10'd                 832;
defparam Ur5_n_13_pp.C8 = 10'd                  51;
defparam Ur5_n_13_pp.C9 = 10'd                 833;
defparam Ur5_n_13_pp.CA = 10'd                   1;
defparam Ur5_n_13_pp.CB = 10'd                 783;
defparam Ur5_n_13_pp.CC = 10'd                 151;
defparam Ur5_n_13_pp.CD = 10'd                 933;
defparam Ur5_n_13_pp.CE = 10'd                 101;
defparam Ur5_n_13_pp.CF = 10'd                 883;
assign lut_val_5_n_13_pp[13] = lut_val_5_n_13_pp[9];
assign lut_val_5_n_13_pp[12] = lut_val_5_n_13_pp[9];
assign lut_val_5_n_13_pp[11] = lut_val_5_n_13_pp[9];
assign lut_val_5_n_13_pp[10] = lut_val_5_n_13_pp[9];
wire [13:0] lut_val_5_n_14_pp;
rom_lut_r_cen Ur5_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[14],sym_res_22_n[14],sym_res_21_n[14],sym_res_20_n[14] } ), .data_out( lut_val_5_n_14_pp[9:0]) ) ;
 defparam Ur5_n_14_pp.DATA_WIDTH = 10;
defparam Ur5_n_14_pp.C0 = 10'd                   0;
defparam Ur5_n_14_pp.C1 = 10'd                 782;
defparam Ur5_n_14_pp.C2 = 10'd                 974;
defparam Ur5_n_14_pp.C3 = 10'd                 732;
defparam Ur5_n_14_pp.C4 = 10'd                 100;
defparam Ur5_n_14_pp.C5 = 10'd                 882;
defparam Ur5_n_14_pp.C6 = 10'd                  50;
defparam Ur5_n_14_pp.C7 = 10'd                 832;
defparam Ur5_n_14_pp.C8 = 10'd                  51;
defparam Ur5_n_14_pp.C9 = 10'd                 833;
defparam Ur5_n_14_pp.CA = 10'd                   1;
defparam Ur5_n_14_pp.CB = 10'd                 783;
defparam Ur5_n_14_pp.CC = 10'd                 151;
defparam Ur5_n_14_pp.CD = 10'd                 933;
defparam Ur5_n_14_pp.CE = 10'd                 101;
defparam Ur5_n_14_pp.CF = 10'd                 883;
assign lut_val_5_n_14_pp[13] = lut_val_5_n_14_pp[9];
assign lut_val_5_n_14_pp[12] = lut_val_5_n_14_pp[9];
assign lut_val_5_n_14_pp[11] = lut_val_5_n_14_pp[9];
assign lut_val_5_n_14_pp[10] = lut_val_5_n_14_pp[9];
wire [13:0] lut_val_5_n_15_pp;
rom_lut_r_cen Ur5_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_23_n[15],sym_res_22_n[15],sym_res_21_n[15],sym_res_20_n[15] } ), .data_out( lut_val_5_n_15_pp[9:0]) ) ;
 defparam Ur5_n_15_pp.DATA_WIDTH = 10;
defparam Ur5_n_15_pp.C0 = 10'd                   0;
defparam Ur5_n_15_pp.C1 = 10'd                 782;
defparam Ur5_n_15_pp.C2 = 10'd                 974;
defparam Ur5_n_15_pp.C3 = 10'd                 732;
defparam Ur5_n_15_pp.C4 = 10'd                 100;
defparam Ur5_n_15_pp.C5 = 10'd                 882;
defparam Ur5_n_15_pp.C6 = 10'd                  50;
defparam Ur5_n_15_pp.C7 = 10'd                 832;
defparam Ur5_n_15_pp.C8 = 10'd                  51;
defparam Ur5_n_15_pp.C9 = 10'd                 833;
defparam Ur5_n_15_pp.CA = 10'd                   1;
defparam Ur5_n_15_pp.CB = 10'd                 783;
defparam Ur5_n_15_pp.CC = 10'd                 151;
defparam Ur5_n_15_pp.CD = 10'd                 933;
defparam Ur5_n_15_pp.CE = 10'd                 101;
defparam Ur5_n_15_pp.CF = 10'd                 883;
assign lut_val_5_n_15_pp[13] = lut_val_5_n_15_pp[9];
assign lut_val_5_n_15_pp[12] = lut_val_5_n_15_pp[9];
assign lut_val_5_n_15_pp[11] = lut_val_5_n_15_pp[9];
assign lut_val_5_n_15_pp[10] = lut_val_5_n_15_pp[9];
wire [13:0] lut_val_6_n_0_pp;
rom_lut_r_cen Ur6_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[0],sym_res_26_n[0],sym_res_25_n[0],sym_res_24_n[0] } ), .data_out( lut_val_6_n_0_pp[10:0]) ) ;
 defparam Ur6_n_0_pp.DATA_WIDTH = 11;
defparam Ur6_n_0_pp.C0 = 11'd                   0;
defparam Ur6_n_0_pp.C1 = 11'd                1941;
defparam Ur6_n_0_pp.C2 = 11'd                1951;
defparam Ur6_n_0_pp.C3 = 11'd                1844;
defparam Ur6_n_0_pp.C4 = 11'd                 216;
defparam Ur6_n_0_pp.C5 = 11'd                 109;
defparam Ur6_n_0_pp.C6 = 11'd                 119;
defparam Ur6_n_0_pp.C7 = 11'd                  12;
defparam Ur6_n_0_pp.C8 = 11'd                 612;
defparam Ur6_n_0_pp.C9 = 11'd                 505;
defparam Ur6_n_0_pp.CA = 11'd                 515;
defparam Ur6_n_0_pp.CB = 11'd                 408;
defparam Ur6_n_0_pp.CC = 11'd                 828;
defparam Ur6_n_0_pp.CD = 11'd                 721;
defparam Ur6_n_0_pp.CE = 11'd                 731;
defparam Ur6_n_0_pp.CF = 11'd                 624;
assign lut_val_6_n_0_pp[13] = lut_val_6_n_0_pp[10];
assign lut_val_6_n_0_pp[12] = lut_val_6_n_0_pp[10];
assign lut_val_6_n_0_pp[11] = lut_val_6_n_0_pp[10];
wire [13:0] lut_val_6_n_1_pp;
rom_lut_r_cen Ur6_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[1],sym_res_26_n[1],sym_res_25_n[1],sym_res_24_n[1] } ), .data_out( lut_val_6_n_1_pp[10:0]) ) ;
 defparam Ur6_n_1_pp.DATA_WIDTH = 11;
defparam Ur6_n_1_pp.C0 = 11'd                   0;
defparam Ur6_n_1_pp.C1 = 11'd                1941;
defparam Ur6_n_1_pp.C2 = 11'd                1951;
defparam Ur6_n_1_pp.C3 = 11'd                1844;
defparam Ur6_n_1_pp.C4 = 11'd                 216;
defparam Ur6_n_1_pp.C5 = 11'd                 109;
defparam Ur6_n_1_pp.C6 = 11'd                 119;
defparam Ur6_n_1_pp.C7 = 11'd                  12;
defparam Ur6_n_1_pp.C8 = 11'd                 612;
defparam Ur6_n_1_pp.C9 = 11'd                 505;
defparam Ur6_n_1_pp.CA = 11'd                 515;
defparam Ur6_n_1_pp.CB = 11'd                 408;
defparam Ur6_n_1_pp.CC = 11'd                 828;
defparam Ur6_n_1_pp.CD = 11'd                 721;
defparam Ur6_n_1_pp.CE = 11'd                 731;
defparam Ur6_n_1_pp.CF = 11'd                 624;
assign lut_val_6_n_1_pp[13] = lut_val_6_n_1_pp[10];
assign lut_val_6_n_1_pp[12] = lut_val_6_n_1_pp[10];
assign lut_val_6_n_1_pp[11] = lut_val_6_n_1_pp[10];
wire [13:0] lut_val_6_n_2_pp;
rom_lut_r_cen Ur6_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[2],sym_res_26_n[2],sym_res_25_n[2],sym_res_24_n[2] } ), .data_out( lut_val_6_n_2_pp[10:0]) ) ;
 defparam Ur6_n_2_pp.DATA_WIDTH = 11;
defparam Ur6_n_2_pp.C0 = 11'd                   0;
defparam Ur6_n_2_pp.C1 = 11'd                1941;
defparam Ur6_n_2_pp.C2 = 11'd                1951;
defparam Ur6_n_2_pp.C3 = 11'd                1844;
defparam Ur6_n_2_pp.C4 = 11'd                 216;
defparam Ur6_n_2_pp.C5 = 11'd                 109;
defparam Ur6_n_2_pp.C6 = 11'd                 119;
defparam Ur6_n_2_pp.C7 = 11'd                  12;
defparam Ur6_n_2_pp.C8 = 11'd                 612;
defparam Ur6_n_2_pp.C9 = 11'd                 505;
defparam Ur6_n_2_pp.CA = 11'd                 515;
defparam Ur6_n_2_pp.CB = 11'd                 408;
defparam Ur6_n_2_pp.CC = 11'd                 828;
defparam Ur6_n_2_pp.CD = 11'd                 721;
defparam Ur6_n_2_pp.CE = 11'd                 731;
defparam Ur6_n_2_pp.CF = 11'd                 624;
assign lut_val_6_n_2_pp[13] = lut_val_6_n_2_pp[10];
assign lut_val_6_n_2_pp[12] = lut_val_6_n_2_pp[10];
assign lut_val_6_n_2_pp[11] = lut_val_6_n_2_pp[10];
wire [13:0] lut_val_6_n_3_pp;
rom_lut_r_cen Ur6_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[3],sym_res_26_n[3],sym_res_25_n[3],sym_res_24_n[3] } ), .data_out( lut_val_6_n_3_pp[10:0]) ) ;
 defparam Ur6_n_3_pp.DATA_WIDTH = 11;
defparam Ur6_n_3_pp.C0 = 11'd                   0;
defparam Ur6_n_3_pp.C1 = 11'd                1941;
defparam Ur6_n_3_pp.C2 = 11'd                1951;
defparam Ur6_n_3_pp.C3 = 11'd                1844;
defparam Ur6_n_3_pp.C4 = 11'd                 216;
defparam Ur6_n_3_pp.C5 = 11'd                 109;
defparam Ur6_n_3_pp.C6 = 11'd                 119;
defparam Ur6_n_3_pp.C7 = 11'd                  12;
defparam Ur6_n_3_pp.C8 = 11'd                 612;
defparam Ur6_n_3_pp.C9 = 11'd                 505;
defparam Ur6_n_3_pp.CA = 11'd                 515;
defparam Ur6_n_3_pp.CB = 11'd                 408;
defparam Ur6_n_3_pp.CC = 11'd                 828;
defparam Ur6_n_3_pp.CD = 11'd                 721;
defparam Ur6_n_3_pp.CE = 11'd                 731;
defparam Ur6_n_3_pp.CF = 11'd                 624;
assign lut_val_6_n_3_pp[13] = lut_val_6_n_3_pp[10];
assign lut_val_6_n_3_pp[12] = lut_val_6_n_3_pp[10];
assign lut_val_6_n_3_pp[11] = lut_val_6_n_3_pp[10];
wire [13:0] lut_val_6_n_4_pp;
rom_lut_r_cen Ur6_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[4],sym_res_26_n[4],sym_res_25_n[4],sym_res_24_n[4] } ), .data_out( lut_val_6_n_4_pp[10:0]) ) ;
 defparam Ur6_n_4_pp.DATA_WIDTH = 11;
defparam Ur6_n_4_pp.C0 = 11'd                   0;
defparam Ur6_n_4_pp.C1 = 11'd                1941;
defparam Ur6_n_4_pp.C2 = 11'd                1951;
defparam Ur6_n_4_pp.C3 = 11'd                1844;
defparam Ur6_n_4_pp.C4 = 11'd                 216;
defparam Ur6_n_4_pp.C5 = 11'd                 109;
defparam Ur6_n_4_pp.C6 = 11'd                 119;
defparam Ur6_n_4_pp.C7 = 11'd                  12;
defparam Ur6_n_4_pp.C8 = 11'd                 612;
defparam Ur6_n_4_pp.C9 = 11'd                 505;
defparam Ur6_n_4_pp.CA = 11'd                 515;
defparam Ur6_n_4_pp.CB = 11'd                 408;
defparam Ur6_n_4_pp.CC = 11'd                 828;
defparam Ur6_n_4_pp.CD = 11'd                 721;
defparam Ur6_n_4_pp.CE = 11'd                 731;
defparam Ur6_n_4_pp.CF = 11'd                 624;
assign lut_val_6_n_4_pp[13] = lut_val_6_n_4_pp[10];
assign lut_val_6_n_4_pp[12] = lut_val_6_n_4_pp[10];
assign lut_val_6_n_4_pp[11] = lut_val_6_n_4_pp[10];
wire [13:0] lut_val_6_n_5_pp;
rom_lut_r_cen Ur6_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[5],sym_res_26_n[5],sym_res_25_n[5],sym_res_24_n[5] } ), .data_out( lut_val_6_n_5_pp[10:0]) ) ;
 defparam Ur6_n_5_pp.DATA_WIDTH = 11;
defparam Ur6_n_5_pp.C0 = 11'd                   0;
defparam Ur6_n_5_pp.C1 = 11'd                1941;
defparam Ur6_n_5_pp.C2 = 11'd                1951;
defparam Ur6_n_5_pp.C3 = 11'd                1844;
defparam Ur6_n_5_pp.C4 = 11'd                 216;
defparam Ur6_n_5_pp.C5 = 11'd                 109;
defparam Ur6_n_5_pp.C6 = 11'd                 119;
defparam Ur6_n_5_pp.C7 = 11'd                  12;
defparam Ur6_n_5_pp.C8 = 11'd                 612;
defparam Ur6_n_5_pp.C9 = 11'd                 505;
defparam Ur6_n_5_pp.CA = 11'd                 515;
defparam Ur6_n_5_pp.CB = 11'd                 408;
defparam Ur6_n_5_pp.CC = 11'd                 828;
defparam Ur6_n_5_pp.CD = 11'd                 721;
defparam Ur6_n_5_pp.CE = 11'd                 731;
defparam Ur6_n_5_pp.CF = 11'd                 624;
assign lut_val_6_n_5_pp[13] = lut_val_6_n_5_pp[10];
assign lut_val_6_n_5_pp[12] = lut_val_6_n_5_pp[10];
assign lut_val_6_n_5_pp[11] = lut_val_6_n_5_pp[10];
wire [13:0] lut_val_6_n_6_pp;
rom_lut_r_cen Ur6_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[6],sym_res_26_n[6],sym_res_25_n[6],sym_res_24_n[6] } ), .data_out( lut_val_6_n_6_pp[10:0]) ) ;
 defparam Ur6_n_6_pp.DATA_WIDTH = 11;
defparam Ur6_n_6_pp.C0 = 11'd                   0;
defparam Ur6_n_6_pp.C1 = 11'd                1941;
defparam Ur6_n_6_pp.C2 = 11'd                1951;
defparam Ur6_n_6_pp.C3 = 11'd                1844;
defparam Ur6_n_6_pp.C4 = 11'd                 216;
defparam Ur6_n_6_pp.C5 = 11'd                 109;
defparam Ur6_n_6_pp.C6 = 11'd                 119;
defparam Ur6_n_6_pp.C7 = 11'd                  12;
defparam Ur6_n_6_pp.C8 = 11'd                 612;
defparam Ur6_n_6_pp.C9 = 11'd                 505;
defparam Ur6_n_6_pp.CA = 11'd                 515;
defparam Ur6_n_6_pp.CB = 11'd                 408;
defparam Ur6_n_6_pp.CC = 11'd                 828;
defparam Ur6_n_6_pp.CD = 11'd                 721;
defparam Ur6_n_6_pp.CE = 11'd                 731;
defparam Ur6_n_6_pp.CF = 11'd                 624;
assign lut_val_6_n_6_pp[13] = lut_val_6_n_6_pp[10];
assign lut_val_6_n_6_pp[12] = lut_val_6_n_6_pp[10];
assign lut_val_6_n_6_pp[11] = lut_val_6_n_6_pp[10];
wire [13:0] lut_val_6_n_7_pp;
rom_lut_r_cen Ur6_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[7],sym_res_26_n[7],sym_res_25_n[7],sym_res_24_n[7] } ), .data_out( lut_val_6_n_7_pp[10:0]) ) ;
 defparam Ur6_n_7_pp.DATA_WIDTH = 11;
defparam Ur6_n_7_pp.C0 = 11'd                   0;
defparam Ur6_n_7_pp.C1 = 11'd                1941;
defparam Ur6_n_7_pp.C2 = 11'd                1951;
defparam Ur6_n_7_pp.C3 = 11'd                1844;
defparam Ur6_n_7_pp.C4 = 11'd                 216;
defparam Ur6_n_7_pp.C5 = 11'd                 109;
defparam Ur6_n_7_pp.C6 = 11'd                 119;
defparam Ur6_n_7_pp.C7 = 11'd                  12;
defparam Ur6_n_7_pp.C8 = 11'd                 612;
defparam Ur6_n_7_pp.C9 = 11'd                 505;
defparam Ur6_n_7_pp.CA = 11'd                 515;
defparam Ur6_n_7_pp.CB = 11'd                 408;
defparam Ur6_n_7_pp.CC = 11'd                 828;
defparam Ur6_n_7_pp.CD = 11'd                 721;
defparam Ur6_n_7_pp.CE = 11'd                 731;
defparam Ur6_n_7_pp.CF = 11'd                 624;
assign lut_val_6_n_7_pp[13] = lut_val_6_n_7_pp[10];
assign lut_val_6_n_7_pp[12] = lut_val_6_n_7_pp[10];
assign lut_val_6_n_7_pp[11] = lut_val_6_n_7_pp[10];
wire [13:0] lut_val_6_n_8_pp;
rom_lut_r_cen Ur6_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[8],sym_res_26_n[8],sym_res_25_n[8],sym_res_24_n[8] } ), .data_out( lut_val_6_n_8_pp[10:0]) ) ;
 defparam Ur6_n_8_pp.DATA_WIDTH = 11;
defparam Ur6_n_8_pp.C0 = 11'd                   0;
defparam Ur6_n_8_pp.C1 = 11'd                1941;
defparam Ur6_n_8_pp.C2 = 11'd                1951;
defparam Ur6_n_8_pp.C3 = 11'd                1844;
defparam Ur6_n_8_pp.C4 = 11'd                 216;
defparam Ur6_n_8_pp.C5 = 11'd                 109;
defparam Ur6_n_8_pp.C6 = 11'd                 119;
defparam Ur6_n_8_pp.C7 = 11'd                  12;
defparam Ur6_n_8_pp.C8 = 11'd                 612;
defparam Ur6_n_8_pp.C9 = 11'd                 505;
defparam Ur6_n_8_pp.CA = 11'd                 515;
defparam Ur6_n_8_pp.CB = 11'd                 408;
defparam Ur6_n_8_pp.CC = 11'd                 828;
defparam Ur6_n_8_pp.CD = 11'd                 721;
defparam Ur6_n_8_pp.CE = 11'd                 731;
defparam Ur6_n_8_pp.CF = 11'd                 624;
assign lut_val_6_n_8_pp[13] = lut_val_6_n_8_pp[10];
assign lut_val_6_n_8_pp[12] = lut_val_6_n_8_pp[10];
assign lut_val_6_n_8_pp[11] = lut_val_6_n_8_pp[10];
wire [13:0] lut_val_6_n_9_pp;
rom_lut_r_cen Ur6_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[9],sym_res_26_n[9],sym_res_25_n[9],sym_res_24_n[9] } ), .data_out( lut_val_6_n_9_pp[10:0]) ) ;
 defparam Ur6_n_9_pp.DATA_WIDTH = 11;
defparam Ur6_n_9_pp.C0 = 11'd                   0;
defparam Ur6_n_9_pp.C1 = 11'd                1941;
defparam Ur6_n_9_pp.C2 = 11'd                1951;
defparam Ur6_n_9_pp.C3 = 11'd                1844;
defparam Ur6_n_9_pp.C4 = 11'd                 216;
defparam Ur6_n_9_pp.C5 = 11'd                 109;
defparam Ur6_n_9_pp.C6 = 11'd                 119;
defparam Ur6_n_9_pp.C7 = 11'd                  12;
defparam Ur6_n_9_pp.C8 = 11'd                 612;
defparam Ur6_n_9_pp.C9 = 11'd                 505;
defparam Ur6_n_9_pp.CA = 11'd                 515;
defparam Ur6_n_9_pp.CB = 11'd                 408;
defparam Ur6_n_9_pp.CC = 11'd                 828;
defparam Ur6_n_9_pp.CD = 11'd                 721;
defparam Ur6_n_9_pp.CE = 11'd                 731;
defparam Ur6_n_9_pp.CF = 11'd                 624;
assign lut_val_6_n_9_pp[13] = lut_val_6_n_9_pp[10];
assign lut_val_6_n_9_pp[12] = lut_val_6_n_9_pp[10];
assign lut_val_6_n_9_pp[11] = lut_val_6_n_9_pp[10];
wire [13:0] lut_val_6_n_10_pp;
rom_lut_r_cen Ur6_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[10],sym_res_26_n[10],sym_res_25_n[10],sym_res_24_n[10] } ), .data_out( lut_val_6_n_10_pp[10:0]) ) ;
 defparam Ur6_n_10_pp.DATA_WIDTH = 11;
defparam Ur6_n_10_pp.C0 = 11'd                   0;
defparam Ur6_n_10_pp.C1 = 11'd                1941;
defparam Ur6_n_10_pp.C2 = 11'd                1951;
defparam Ur6_n_10_pp.C3 = 11'd                1844;
defparam Ur6_n_10_pp.C4 = 11'd                 216;
defparam Ur6_n_10_pp.C5 = 11'd                 109;
defparam Ur6_n_10_pp.C6 = 11'd                 119;
defparam Ur6_n_10_pp.C7 = 11'd                  12;
defparam Ur6_n_10_pp.C8 = 11'd                 612;
defparam Ur6_n_10_pp.C9 = 11'd                 505;
defparam Ur6_n_10_pp.CA = 11'd                 515;
defparam Ur6_n_10_pp.CB = 11'd                 408;
defparam Ur6_n_10_pp.CC = 11'd                 828;
defparam Ur6_n_10_pp.CD = 11'd                 721;
defparam Ur6_n_10_pp.CE = 11'd                 731;
defparam Ur6_n_10_pp.CF = 11'd                 624;
assign lut_val_6_n_10_pp[13] = lut_val_6_n_10_pp[10];
assign lut_val_6_n_10_pp[12] = lut_val_6_n_10_pp[10];
assign lut_val_6_n_10_pp[11] = lut_val_6_n_10_pp[10];
wire [13:0] lut_val_6_n_11_pp;
rom_lut_r_cen Ur6_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[11],sym_res_26_n[11],sym_res_25_n[11],sym_res_24_n[11] } ), .data_out( lut_val_6_n_11_pp[10:0]) ) ;
 defparam Ur6_n_11_pp.DATA_WIDTH = 11;
defparam Ur6_n_11_pp.C0 = 11'd                   0;
defparam Ur6_n_11_pp.C1 = 11'd                1941;
defparam Ur6_n_11_pp.C2 = 11'd                1951;
defparam Ur6_n_11_pp.C3 = 11'd                1844;
defparam Ur6_n_11_pp.C4 = 11'd                 216;
defparam Ur6_n_11_pp.C5 = 11'd                 109;
defparam Ur6_n_11_pp.C6 = 11'd                 119;
defparam Ur6_n_11_pp.C7 = 11'd                  12;
defparam Ur6_n_11_pp.C8 = 11'd                 612;
defparam Ur6_n_11_pp.C9 = 11'd                 505;
defparam Ur6_n_11_pp.CA = 11'd                 515;
defparam Ur6_n_11_pp.CB = 11'd                 408;
defparam Ur6_n_11_pp.CC = 11'd                 828;
defparam Ur6_n_11_pp.CD = 11'd                 721;
defparam Ur6_n_11_pp.CE = 11'd                 731;
defparam Ur6_n_11_pp.CF = 11'd                 624;
assign lut_val_6_n_11_pp[13] = lut_val_6_n_11_pp[10];
assign lut_val_6_n_11_pp[12] = lut_val_6_n_11_pp[10];
assign lut_val_6_n_11_pp[11] = lut_val_6_n_11_pp[10];
wire [13:0] lut_val_6_n_12_pp;
rom_lut_r_cen Ur6_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[12],sym_res_26_n[12],sym_res_25_n[12],sym_res_24_n[12] } ), .data_out( lut_val_6_n_12_pp[10:0]) ) ;
 defparam Ur6_n_12_pp.DATA_WIDTH = 11;
defparam Ur6_n_12_pp.C0 = 11'd                   0;
defparam Ur6_n_12_pp.C1 = 11'd                1941;
defparam Ur6_n_12_pp.C2 = 11'd                1951;
defparam Ur6_n_12_pp.C3 = 11'd                1844;
defparam Ur6_n_12_pp.C4 = 11'd                 216;
defparam Ur6_n_12_pp.C5 = 11'd                 109;
defparam Ur6_n_12_pp.C6 = 11'd                 119;
defparam Ur6_n_12_pp.C7 = 11'd                  12;
defparam Ur6_n_12_pp.C8 = 11'd                 612;
defparam Ur6_n_12_pp.C9 = 11'd                 505;
defparam Ur6_n_12_pp.CA = 11'd                 515;
defparam Ur6_n_12_pp.CB = 11'd                 408;
defparam Ur6_n_12_pp.CC = 11'd                 828;
defparam Ur6_n_12_pp.CD = 11'd                 721;
defparam Ur6_n_12_pp.CE = 11'd                 731;
defparam Ur6_n_12_pp.CF = 11'd                 624;
assign lut_val_6_n_12_pp[13] = lut_val_6_n_12_pp[10];
assign lut_val_6_n_12_pp[12] = lut_val_6_n_12_pp[10];
assign lut_val_6_n_12_pp[11] = lut_val_6_n_12_pp[10];
wire [13:0] lut_val_6_n_13_pp;
rom_lut_r_cen Ur6_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[13],sym_res_26_n[13],sym_res_25_n[13],sym_res_24_n[13] } ), .data_out( lut_val_6_n_13_pp[10:0]) ) ;
 defparam Ur6_n_13_pp.DATA_WIDTH = 11;
defparam Ur6_n_13_pp.C0 = 11'd                   0;
defparam Ur6_n_13_pp.C1 = 11'd                1941;
defparam Ur6_n_13_pp.C2 = 11'd                1951;
defparam Ur6_n_13_pp.C3 = 11'd                1844;
defparam Ur6_n_13_pp.C4 = 11'd                 216;
defparam Ur6_n_13_pp.C5 = 11'd                 109;
defparam Ur6_n_13_pp.C6 = 11'd                 119;
defparam Ur6_n_13_pp.C7 = 11'd                  12;
defparam Ur6_n_13_pp.C8 = 11'd                 612;
defparam Ur6_n_13_pp.C9 = 11'd                 505;
defparam Ur6_n_13_pp.CA = 11'd                 515;
defparam Ur6_n_13_pp.CB = 11'd                 408;
defparam Ur6_n_13_pp.CC = 11'd                 828;
defparam Ur6_n_13_pp.CD = 11'd                 721;
defparam Ur6_n_13_pp.CE = 11'd                 731;
defparam Ur6_n_13_pp.CF = 11'd                 624;
assign lut_val_6_n_13_pp[13] = lut_val_6_n_13_pp[10];
assign lut_val_6_n_13_pp[12] = lut_val_6_n_13_pp[10];
assign lut_val_6_n_13_pp[11] = lut_val_6_n_13_pp[10];
wire [13:0] lut_val_6_n_14_pp;
rom_lut_r_cen Ur6_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[14],sym_res_26_n[14],sym_res_25_n[14],sym_res_24_n[14] } ), .data_out( lut_val_6_n_14_pp[10:0]) ) ;
 defparam Ur6_n_14_pp.DATA_WIDTH = 11;
defparam Ur6_n_14_pp.C0 = 11'd                   0;
defparam Ur6_n_14_pp.C1 = 11'd                1941;
defparam Ur6_n_14_pp.C2 = 11'd                1951;
defparam Ur6_n_14_pp.C3 = 11'd                1844;
defparam Ur6_n_14_pp.C4 = 11'd                 216;
defparam Ur6_n_14_pp.C5 = 11'd                 109;
defparam Ur6_n_14_pp.C6 = 11'd                 119;
defparam Ur6_n_14_pp.C7 = 11'd                  12;
defparam Ur6_n_14_pp.C8 = 11'd                 612;
defparam Ur6_n_14_pp.C9 = 11'd                 505;
defparam Ur6_n_14_pp.CA = 11'd                 515;
defparam Ur6_n_14_pp.CB = 11'd                 408;
defparam Ur6_n_14_pp.CC = 11'd                 828;
defparam Ur6_n_14_pp.CD = 11'd                 721;
defparam Ur6_n_14_pp.CE = 11'd                 731;
defparam Ur6_n_14_pp.CF = 11'd                 624;
assign lut_val_6_n_14_pp[13] = lut_val_6_n_14_pp[10];
assign lut_val_6_n_14_pp[12] = lut_val_6_n_14_pp[10];
assign lut_val_6_n_14_pp[11] = lut_val_6_n_14_pp[10];
wire [13:0] lut_val_6_n_15_pp;
rom_lut_r_cen Ur6_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_27_n[15],sym_res_26_n[15],sym_res_25_n[15],sym_res_24_n[15] } ), .data_out( lut_val_6_n_15_pp[10:0]) ) ;
 defparam Ur6_n_15_pp.DATA_WIDTH = 11;
defparam Ur6_n_15_pp.C0 = 11'd                   0;
defparam Ur6_n_15_pp.C1 = 11'd                1941;
defparam Ur6_n_15_pp.C2 = 11'd                1951;
defparam Ur6_n_15_pp.C3 = 11'd                1844;
defparam Ur6_n_15_pp.C4 = 11'd                 216;
defparam Ur6_n_15_pp.C5 = 11'd                 109;
defparam Ur6_n_15_pp.C6 = 11'd                 119;
defparam Ur6_n_15_pp.C7 = 11'd                  12;
defparam Ur6_n_15_pp.C8 = 11'd                 612;
defparam Ur6_n_15_pp.C9 = 11'd                 505;
defparam Ur6_n_15_pp.CA = 11'd                 515;
defparam Ur6_n_15_pp.CB = 11'd                 408;
defparam Ur6_n_15_pp.CC = 11'd                 828;
defparam Ur6_n_15_pp.CD = 11'd                 721;
defparam Ur6_n_15_pp.CE = 11'd                 731;
defparam Ur6_n_15_pp.CF = 11'd                 624;
assign lut_val_6_n_15_pp[13] = lut_val_6_n_15_pp[10];
assign lut_val_6_n_15_pp[12] = lut_val_6_n_15_pp[10];
assign lut_val_6_n_15_pp[11] = lut_val_6_n_15_pp[10];
wire [13:0] lut_val_7_n_0_pp;
rom_lut_r_cen Ur7_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[0],sym_res_30_n[0],sym_res_29_n[0],sym_res_28_n[0] } ), .data_out( lut_val_7_n_0_pp[10:0]) ) ;
 defparam Ur7_n_0_pp.DATA_WIDTH = 11;
defparam Ur7_n_0_pp.C0 = 11'd                   0;
defparam Ur7_n_0_pp.C1 = 11'd                 684;
defparam Ur7_n_0_pp.C2 = 11'd                 302;
defparam Ur7_n_0_pp.C3 = 11'd                 986;
defparam Ur7_n_0_pp.C4 = 11'd                1876;
defparam Ur7_n_0_pp.C5 = 11'd                 512;
defparam Ur7_n_0_pp.C6 = 11'd                 130;
defparam Ur7_n_0_pp.C7 = 11'd                 814;
defparam Ur7_n_0_pp.C8 = 11'd                1814;
defparam Ur7_n_0_pp.C9 = 11'd                 450;
defparam Ur7_n_0_pp.CA = 11'd                  68;
defparam Ur7_n_0_pp.CB = 11'd                 752;
defparam Ur7_n_0_pp.CC = 11'd                1642;
defparam Ur7_n_0_pp.CD = 11'd                 278;
defparam Ur7_n_0_pp.CE = 11'd                1944;
defparam Ur7_n_0_pp.CF = 11'd                 580;
assign lut_val_7_n_0_pp[13] = lut_val_7_n_0_pp[10];
assign lut_val_7_n_0_pp[12] = lut_val_7_n_0_pp[10];
assign lut_val_7_n_0_pp[11] = lut_val_7_n_0_pp[10];
wire [13:0] lut_val_7_n_1_pp;
rom_lut_r_cen Ur7_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[1],sym_res_30_n[1],sym_res_29_n[1],sym_res_28_n[1] } ), .data_out( lut_val_7_n_1_pp[10:0]) ) ;
 defparam Ur7_n_1_pp.DATA_WIDTH = 11;
defparam Ur7_n_1_pp.C0 = 11'd                   0;
defparam Ur7_n_1_pp.C1 = 11'd                 684;
defparam Ur7_n_1_pp.C2 = 11'd                 302;
defparam Ur7_n_1_pp.C3 = 11'd                 986;
defparam Ur7_n_1_pp.C4 = 11'd                1876;
defparam Ur7_n_1_pp.C5 = 11'd                 512;
defparam Ur7_n_1_pp.C6 = 11'd                 130;
defparam Ur7_n_1_pp.C7 = 11'd                 814;
defparam Ur7_n_1_pp.C8 = 11'd                1814;
defparam Ur7_n_1_pp.C9 = 11'd                 450;
defparam Ur7_n_1_pp.CA = 11'd                  68;
defparam Ur7_n_1_pp.CB = 11'd                 752;
defparam Ur7_n_1_pp.CC = 11'd                1642;
defparam Ur7_n_1_pp.CD = 11'd                 278;
defparam Ur7_n_1_pp.CE = 11'd                1944;
defparam Ur7_n_1_pp.CF = 11'd                 580;
assign lut_val_7_n_1_pp[13] = lut_val_7_n_1_pp[10];
assign lut_val_7_n_1_pp[12] = lut_val_7_n_1_pp[10];
assign lut_val_7_n_1_pp[11] = lut_val_7_n_1_pp[10];
wire [13:0] lut_val_7_n_2_pp;
rom_lut_r_cen Ur7_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[2],sym_res_30_n[2],sym_res_29_n[2],sym_res_28_n[2] } ), .data_out( lut_val_7_n_2_pp[10:0]) ) ;
 defparam Ur7_n_2_pp.DATA_WIDTH = 11;
defparam Ur7_n_2_pp.C0 = 11'd                   0;
defparam Ur7_n_2_pp.C1 = 11'd                 684;
defparam Ur7_n_2_pp.C2 = 11'd                 302;
defparam Ur7_n_2_pp.C3 = 11'd                 986;
defparam Ur7_n_2_pp.C4 = 11'd                1876;
defparam Ur7_n_2_pp.C5 = 11'd                 512;
defparam Ur7_n_2_pp.C6 = 11'd                 130;
defparam Ur7_n_2_pp.C7 = 11'd                 814;
defparam Ur7_n_2_pp.C8 = 11'd                1814;
defparam Ur7_n_2_pp.C9 = 11'd                 450;
defparam Ur7_n_2_pp.CA = 11'd                  68;
defparam Ur7_n_2_pp.CB = 11'd                 752;
defparam Ur7_n_2_pp.CC = 11'd                1642;
defparam Ur7_n_2_pp.CD = 11'd                 278;
defparam Ur7_n_2_pp.CE = 11'd                1944;
defparam Ur7_n_2_pp.CF = 11'd                 580;
assign lut_val_7_n_2_pp[13] = lut_val_7_n_2_pp[10];
assign lut_val_7_n_2_pp[12] = lut_val_7_n_2_pp[10];
assign lut_val_7_n_2_pp[11] = lut_val_7_n_2_pp[10];
wire [13:0] lut_val_7_n_3_pp;
rom_lut_r_cen Ur7_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[3],sym_res_30_n[3],sym_res_29_n[3],sym_res_28_n[3] } ), .data_out( lut_val_7_n_3_pp[10:0]) ) ;
 defparam Ur7_n_3_pp.DATA_WIDTH = 11;
defparam Ur7_n_3_pp.C0 = 11'd                   0;
defparam Ur7_n_3_pp.C1 = 11'd                 684;
defparam Ur7_n_3_pp.C2 = 11'd                 302;
defparam Ur7_n_3_pp.C3 = 11'd                 986;
defparam Ur7_n_3_pp.C4 = 11'd                1876;
defparam Ur7_n_3_pp.C5 = 11'd                 512;
defparam Ur7_n_3_pp.C6 = 11'd                 130;
defparam Ur7_n_3_pp.C7 = 11'd                 814;
defparam Ur7_n_3_pp.C8 = 11'd                1814;
defparam Ur7_n_3_pp.C9 = 11'd                 450;
defparam Ur7_n_3_pp.CA = 11'd                  68;
defparam Ur7_n_3_pp.CB = 11'd                 752;
defparam Ur7_n_3_pp.CC = 11'd                1642;
defparam Ur7_n_3_pp.CD = 11'd                 278;
defparam Ur7_n_3_pp.CE = 11'd                1944;
defparam Ur7_n_3_pp.CF = 11'd                 580;
assign lut_val_7_n_3_pp[13] = lut_val_7_n_3_pp[10];
assign lut_val_7_n_3_pp[12] = lut_val_7_n_3_pp[10];
assign lut_val_7_n_3_pp[11] = lut_val_7_n_3_pp[10];
wire [13:0] lut_val_7_n_4_pp;
rom_lut_r_cen Ur7_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[4],sym_res_30_n[4],sym_res_29_n[4],sym_res_28_n[4] } ), .data_out( lut_val_7_n_4_pp[10:0]) ) ;
 defparam Ur7_n_4_pp.DATA_WIDTH = 11;
defparam Ur7_n_4_pp.C0 = 11'd                   0;
defparam Ur7_n_4_pp.C1 = 11'd                 684;
defparam Ur7_n_4_pp.C2 = 11'd                 302;
defparam Ur7_n_4_pp.C3 = 11'd                 986;
defparam Ur7_n_4_pp.C4 = 11'd                1876;
defparam Ur7_n_4_pp.C5 = 11'd                 512;
defparam Ur7_n_4_pp.C6 = 11'd                 130;
defparam Ur7_n_4_pp.C7 = 11'd                 814;
defparam Ur7_n_4_pp.C8 = 11'd                1814;
defparam Ur7_n_4_pp.C9 = 11'd                 450;
defparam Ur7_n_4_pp.CA = 11'd                  68;
defparam Ur7_n_4_pp.CB = 11'd                 752;
defparam Ur7_n_4_pp.CC = 11'd                1642;
defparam Ur7_n_4_pp.CD = 11'd                 278;
defparam Ur7_n_4_pp.CE = 11'd                1944;
defparam Ur7_n_4_pp.CF = 11'd                 580;
assign lut_val_7_n_4_pp[13] = lut_val_7_n_4_pp[10];
assign lut_val_7_n_4_pp[12] = lut_val_7_n_4_pp[10];
assign lut_val_7_n_4_pp[11] = lut_val_7_n_4_pp[10];
wire [13:0] lut_val_7_n_5_pp;
rom_lut_r_cen Ur7_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[5],sym_res_30_n[5],sym_res_29_n[5],sym_res_28_n[5] } ), .data_out( lut_val_7_n_5_pp[10:0]) ) ;
 defparam Ur7_n_5_pp.DATA_WIDTH = 11;
defparam Ur7_n_5_pp.C0 = 11'd                   0;
defparam Ur7_n_5_pp.C1 = 11'd                 684;
defparam Ur7_n_5_pp.C2 = 11'd                 302;
defparam Ur7_n_5_pp.C3 = 11'd                 986;
defparam Ur7_n_5_pp.C4 = 11'd                1876;
defparam Ur7_n_5_pp.C5 = 11'd                 512;
defparam Ur7_n_5_pp.C6 = 11'd                 130;
defparam Ur7_n_5_pp.C7 = 11'd                 814;
defparam Ur7_n_5_pp.C8 = 11'd                1814;
defparam Ur7_n_5_pp.C9 = 11'd                 450;
defparam Ur7_n_5_pp.CA = 11'd                  68;
defparam Ur7_n_5_pp.CB = 11'd                 752;
defparam Ur7_n_5_pp.CC = 11'd                1642;
defparam Ur7_n_5_pp.CD = 11'd                 278;
defparam Ur7_n_5_pp.CE = 11'd                1944;
defparam Ur7_n_5_pp.CF = 11'd                 580;
assign lut_val_7_n_5_pp[13] = lut_val_7_n_5_pp[10];
assign lut_val_7_n_5_pp[12] = lut_val_7_n_5_pp[10];
assign lut_val_7_n_5_pp[11] = lut_val_7_n_5_pp[10];
wire [13:0] lut_val_7_n_6_pp;
rom_lut_r_cen Ur7_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[6],sym_res_30_n[6],sym_res_29_n[6],sym_res_28_n[6] } ), .data_out( lut_val_7_n_6_pp[10:0]) ) ;
 defparam Ur7_n_6_pp.DATA_WIDTH = 11;
defparam Ur7_n_6_pp.C0 = 11'd                   0;
defparam Ur7_n_6_pp.C1 = 11'd                 684;
defparam Ur7_n_6_pp.C2 = 11'd                 302;
defparam Ur7_n_6_pp.C3 = 11'd                 986;
defparam Ur7_n_6_pp.C4 = 11'd                1876;
defparam Ur7_n_6_pp.C5 = 11'd                 512;
defparam Ur7_n_6_pp.C6 = 11'd                 130;
defparam Ur7_n_6_pp.C7 = 11'd                 814;
defparam Ur7_n_6_pp.C8 = 11'd                1814;
defparam Ur7_n_6_pp.C9 = 11'd                 450;
defparam Ur7_n_6_pp.CA = 11'd                  68;
defparam Ur7_n_6_pp.CB = 11'd                 752;
defparam Ur7_n_6_pp.CC = 11'd                1642;
defparam Ur7_n_6_pp.CD = 11'd                 278;
defparam Ur7_n_6_pp.CE = 11'd                1944;
defparam Ur7_n_6_pp.CF = 11'd                 580;
assign lut_val_7_n_6_pp[13] = lut_val_7_n_6_pp[10];
assign lut_val_7_n_6_pp[12] = lut_val_7_n_6_pp[10];
assign lut_val_7_n_6_pp[11] = lut_val_7_n_6_pp[10];
wire [13:0] lut_val_7_n_7_pp;
rom_lut_r_cen Ur7_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[7],sym_res_30_n[7],sym_res_29_n[7],sym_res_28_n[7] } ), .data_out( lut_val_7_n_7_pp[10:0]) ) ;
 defparam Ur7_n_7_pp.DATA_WIDTH = 11;
defparam Ur7_n_7_pp.C0 = 11'd                   0;
defparam Ur7_n_7_pp.C1 = 11'd                 684;
defparam Ur7_n_7_pp.C2 = 11'd                 302;
defparam Ur7_n_7_pp.C3 = 11'd                 986;
defparam Ur7_n_7_pp.C4 = 11'd                1876;
defparam Ur7_n_7_pp.C5 = 11'd                 512;
defparam Ur7_n_7_pp.C6 = 11'd                 130;
defparam Ur7_n_7_pp.C7 = 11'd                 814;
defparam Ur7_n_7_pp.C8 = 11'd                1814;
defparam Ur7_n_7_pp.C9 = 11'd                 450;
defparam Ur7_n_7_pp.CA = 11'd                  68;
defparam Ur7_n_7_pp.CB = 11'd                 752;
defparam Ur7_n_7_pp.CC = 11'd                1642;
defparam Ur7_n_7_pp.CD = 11'd                 278;
defparam Ur7_n_7_pp.CE = 11'd                1944;
defparam Ur7_n_7_pp.CF = 11'd                 580;
assign lut_val_7_n_7_pp[13] = lut_val_7_n_7_pp[10];
assign lut_val_7_n_7_pp[12] = lut_val_7_n_7_pp[10];
assign lut_val_7_n_7_pp[11] = lut_val_7_n_7_pp[10];
wire [13:0] lut_val_7_n_8_pp;
rom_lut_r_cen Ur7_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[8],sym_res_30_n[8],sym_res_29_n[8],sym_res_28_n[8] } ), .data_out( lut_val_7_n_8_pp[10:0]) ) ;
 defparam Ur7_n_8_pp.DATA_WIDTH = 11;
defparam Ur7_n_8_pp.C0 = 11'd                   0;
defparam Ur7_n_8_pp.C1 = 11'd                 684;
defparam Ur7_n_8_pp.C2 = 11'd                 302;
defparam Ur7_n_8_pp.C3 = 11'd                 986;
defparam Ur7_n_8_pp.C4 = 11'd                1876;
defparam Ur7_n_8_pp.C5 = 11'd                 512;
defparam Ur7_n_8_pp.C6 = 11'd                 130;
defparam Ur7_n_8_pp.C7 = 11'd                 814;
defparam Ur7_n_8_pp.C8 = 11'd                1814;
defparam Ur7_n_8_pp.C9 = 11'd                 450;
defparam Ur7_n_8_pp.CA = 11'd                  68;
defparam Ur7_n_8_pp.CB = 11'd                 752;
defparam Ur7_n_8_pp.CC = 11'd                1642;
defparam Ur7_n_8_pp.CD = 11'd                 278;
defparam Ur7_n_8_pp.CE = 11'd                1944;
defparam Ur7_n_8_pp.CF = 11'd                 580;
assign lut_val_7_n_8_pp[13] = lut_val_7_n_8_pp[10];
assign lut_val_7_n_8_pp[12] = lut_val_7_n_8_pp[10];
assign lut_val_7_n_8_pp[11] = lut_val_7_n_8_pp[10];
wire [13:0] lut_val_7_n_9_pp;
rom_lut_r_cen Ur7_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[9],sym_res_30_n[9],sym_res_29_n[9],sym_res_28_n[9] } ), .data_out( lut_val_7_n_9_pp[10:0]) ) ;
 defparam Ur7_n_9_pp.DATA_WIDTH = 11;
defparam Ur7_n_9_pp.C0 = 11'd                   0;
defparam Ur7_n_9_pp.C1 = 11'd                 684;
defparam Ur7_n_9_pp.C2 = 11'd                 302;
defparam Ur7_n_9_pp.C3 = 11'd                 986;
defparam Ur7_n_9_pp.C4 = 11'd                1876;
defparam Ur7_n_9_pp.C5 = 11'd                 512;
defparam Ur7_n_9_pp.C6 = 11'd                 130;
defparam Ur7_n_9_pp.C7 = 11'd                 814;
defparam Ur7_n_9_pp.C8 = 11'd                1814;
defparam Ur7_n_9_pp.C9 = 11'd                 450;
defparam Ur7_n_9_pp.CA = 11'd                  68;
defparam Ur7_n_9_pp.CB = 11'd                 752;
defparam Ur7_n_9_pp.CC = 11'd                1642;
defparam Ur7_n_9_pp.CD = 11'd                 278;
defparam Ur7_n_9_pp.CE = 11'd                1944;
defparam Ur7_n_9_pp.CF = 11'd                 580;
assign lut_val_7_n_9_pp[13] = lut_val_7_n_9_pp[10];
assign lut_val_7_n_9_pp[12] = lut_val_7_n_9_pp[10];
assign lut_val_7_n_9_pp[11] = lut_val_7_n_9_pp[10];
wire [13:0] lut_val_7_n_10_pp;
rom_lut_r_cen Ur7_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[10],sym_res_30_n[10],sym_res_29_n[10],sym_res_28_n[10] } ), .data_out( lut_val_7_n_10_pp[10:0]) ) ;
 defparam Ur7_n_10_pp.DATA_WIDTH = 11;
defparam Ur7_n_10_pp.C0 = 11'd                   0;
defparam Ur7_n_10_pp.C1 = 11'd                 684;
defparam Ur7_n_10_pp.C2 = 11'd                 302;
defparam Ur7_n_10_pp.C3 = 11'd                 986;
defparam Ur7_n_10_pp.C4 = 11'd                1876;
defparam Ur7_n_10_pp.C5 = 11'd                 512;
defparam Ur7_n_10_pp.C6 = 11'd                 130;
defparam Ur7_n_10_pp.C7 = 11'd                 814;
defparam Ur7_n_10_pp.C8 = 11'd                1814;
defparam Ur7_n_10_pp.C9 = 11'd                 450;
defparam Ur7_n_10_pp.CA = 11'd                  68;
defparam Ur7_n_10_pp.CB = 11'd                 752;
defparam Ur7_n_10_pp.CC = 11'd                1642;
defparam Ur7_n_10_pp.CD = 11'd                 278;
defparam Ur7_n_10_pp.CE = 11'd                1944;
defparam Ur7_n_10_pp.CF = 11'd                 580;
assign lut_val_7_n_10_pp[13] = lut_val_7_n_10_pp[10];
assign lut_val_7_n_10_pp[12] = lut_val_7_n_10_pp[10];
assign lut_val_7_n_10_pp[11] = lut_val_7_n_10_pp[10];
wire [13:0] lut_val_7_n_11_pp;
rom_lut_r_cen Ur7_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[11],sym_res_30_n[11],sym_res_29_n[11],sym_res_28_n[11] } ), .data_out( lut_val_7_n_11_pp[10:0]) ) ;
 defparam Ur7_n_11_pp.DATA_WIDTH = 11;
defparam Ur7_n_11_pp.C0 = 11'd                   0;
defparam Ur7_n_11_pp.C1 = 11'd                 684;
defparam Ur7_n_11_pp.C2 = 11'd                 302;
defparam Ur7_n_11_pp.C3 = 11'd                 986;
defparam Ur7_n_11_pp.C4 = 11'd                1876;
defparam Ur7_n_11_pp.C5 = 11'd                 512;
defparam Ur7_n_11_pp.C6 = 11'd                 130;
defparam Ur7_n_11_pp.C7 = 11'd                 814;
defparam Ur7_n_11_pp.C8 = 11'd                1814;
defparam Ur7_n_11_pp.C9 = 11'd                 450;
defparam Ur7_n_11_pp.CA = 11'd                  68;
defparam Ur7_n_11_pp.CB = 11'd                 752;
defparam Ur7_n_11_pp.CC = 11'd                1642;
defparam Ur7_n_11_pp.CD = 11'd                 278;
defparam Ur7_n_11_pp.CE = 11'd                1944;
defparam Ur7_n_11_pp.CF = 11'd                 580;
assign lut_val_7_n_11_pp[13] = lut_val_7_n_11_pp[10];
assign lut_val_7_n_11_pp[12] = lut_val_7_n_11_pp[10];
assign lut_val_7_n_11_pp[11] = lut_val_7_n_11_pp[10];
wire [13:0] lut_val_7_n_12_pp;
rom_lut_r_cen Ur7_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[12],sym_res_30_n[12],sym_res_29_n[12],sym_res_28_n[12] } ), .data_out( lut_val_7_n_12_pp[10:0]) ) ;
 defparam Ur7_n_12_pp.DATA_WIDTH = 11;
defparam Ur7_n_12_pp.C0 = 11'd                   0;
defparam Ur7_n_12_pp.C1 = 11'd                 684;
defparam Ur7_n_12_pp.C2 = 11'd                 302;
defparam Ur7_n_12_pp.C3 = 11'd                 986;
defparam Ur7_n_12_pp.C4 = 11'd                1876;
defparam Ur7_n_12_pp.C5 = 11'd                 512;
defparam Ur7_n_12_pp.C6 = 11'd                 130;
defparam Ur7_n_12_pp.C7 = 11'd                 814;
defparam Ur7_n_12_pp.C8 = 11'd                1814;
defparam Ur7_n_12_pp.C9 = 11'd                 450;
defparam Ur7_n_12_pp.CA = 11'd                  68;
defparam Ur7_n_12_pp.CB = 11'd                 752;
defparam Ur7_n_12_pp.CC = 11'd                1642;
defparam Ur7_n_12_pp.CD = 11'd                 278;
defparam Ur7_n_12_pp.CE = 11'd                1944;
defparam Ur7_n_12_pp.CF = 11'd                 580;
assign lut_val_7_n_12_pp[13] = lut_val_7_n_12_pp[10];
assign lut_val_7_n_12_pp[12] = lut_val_7_n_12_pp[10];
assign lut_val_7_n_12_pp[11] = lut_val_7_n_12_pp[10];
wire [13:0] lut_val_7_n_13_pp;
rom_lut_r_cen Ur7_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[13],sym_res_30_n[13],sym_res_29_n[13],sym_res_28_n[13] } ), .data_out( lut_val_7_n_13_pp[10:0]) ) ;
 defparam Ur7_n_13_pp.DATA_WIDTH = 11;
defparam Ur7_n_13_pp.C0 = 11'd                   0;
defparam Ur7_n_13_pp.C1 = 11'd                 684;
defparam Ur7_n_13_pp.C2 = 11'd                 302;
defparam Ur7_n_13_pp.C3 = 11'd                 986;
defparam Ur7_n_13_pp.C4 = 11'd                1876;
defparam Ur7_n_13_pp.C5 = 11'd                 512;
defparam Ur7_n_13_pp.C6 = 11'd                 130;
defparam Ur7_n_13_pp.C7 = 11'd                 814;
defparam Ur7_n_13_pp.C8 = 11'd                1814;
defparam Ur7_n_13_pp.C9 = 11'd                 450;
defparam Ur7_n_13_pp.CA = 11'd                  68;
defparam Ur7_n_13_pp.CB = 11'd                 752;
defparam Ur7_n_13_pp.CC = 11'd                1642;
defparam Ur7_n_13_pp.CD = 11'd                 278;
defparam Ur7_n_13_pp.CE = 11'd                1944;
defparam Ur7_n_13_pp.CF = 11'd                 580;
assign lut_val_7_n_13_pp[13] = lut_val_7_n_13_pp[10];
assign lut_val_7_n_13_pp[12] = lut_val_7_n_13_pp[10];
assign lut_val_7_n_13_pp[11] = lut_val_7_n_13_pp[10];
wire [13:0] lut_val_7_n_14_pp;
rom_lut_r_cen Ur7_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[14],sym_res_30_n[14],sym_res_29_n[14],sym_res_28_n[14] } ), .data_out( lut_val_7_n_14_pp[10:0]) ) ;
 defparam Ur7_n_14_pp.DATA_WIDTH = 11;
defparam Ur7_n_14_pp.C0 = 11'd                   0;
defparam Ur7_n_14_pp.C1 = 11'd                 684;
defparam Ur7_n_14_pp.C2 = 11'd                 302;
defparam Ur7_n_14_pp.C3 = 11'd                 986;
defparam Ur7_n_14_pp.C4 = 11'd                1876;
defparam Ur7_n_14_pp.C5 = 11'd                 512;
defparam Ur7_n_14_pp.C6 = 11'd                 130;
defparam Ur7_n_14_pp.C7 = 11'd                 814;
defparam Ur7_n_14_pp.C8 = 11'd                1814;
defparam Ur7_n_14_pp.C9 = 11'd                 450;
defparam Ur7_n_14_pp.CA = 11'd                  68;
defparam Ur7_n_14_pp.CB = 11'd                 752;
defparam Ur7_n_14_pp.CC = 11'd                1642;
defparam Ur7_n_14_pp.CD = 11'd                 278;
defparam Ur7_n_14_pp.CE = 11'd                1944;
defparam Ur7_n_14_pp.CF = 11'd                 580;
assign lut_val_7_n_14_pp[13] = lut_val_7_n_14_pp[10];
assign lut_val_7_n_14_pp[12] = lut_val_7_n_14_pp[10];
assign lut_val_7_n_14_pp[11] = lut_val_7_n_14_pp[10];
wire [13:0] lut_val_7_n_15_pp;
rom_lut_r_cen Ur7_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_31_n[15],sym_res_30_n[15],sym_res_29_n[15],sym_res_28_n[15] } ), .data_out( lut_val_7_n_15_pp[10:0]) ) ;
 defparam Ur7_n_15_pp.DATA_WIDTH = 11;
defparam Ur7_n_15_pp.C0 = 11'd                   0;
defparam Ur7_n_15_pp.C1 = 11'd                 684;
defparam Ur7_n_15_pp.C2 = 11'd                 302;
defparam Ur7_n_15_pp.C3 = 11'd                 986;
defparam Ur7_n_15_pp.C4 = 11'd                1876;
defparam Ur7_n_15_pp.C5 = 11'd                 512;
defparam Ur7_n_15_pp.C6 = 11'd                 130;
defparam Ur7_n_15_pp.C7 = 11'd                 814;
defparam Ur7_n_15_pp.C8 = 11'd                1814;
defparam Ur7_n_15_pp.C9 = 11'd                 450;
defparam Ur7_n_15_pp.CA = 11'd                  68;
defparam Ur7_n_15_pp.CB = 11'd                 752;
defparam Ur7_n_15_pp.CC = 11'd                1642;
defparam Ur7_n_15_pp.CD = 11'd                 278;
defparam Ur7_n_15_pp.CE = 11'd                1944;
defparam Ur7_n_15_pp.CF = 11'd                 580;
assign lut_val_7_n_15_pp[13] = lut_val_7_n_15_pp[10];
assign lut_val_7_n_15_pp[12] = lut_val_7_n_15_pp[10];
assign lut_val_7_n_15_pp[11] = lut_val_7_n_15_pp[10];
wire [13:0] lut_val_8_n_0_pp;
rom_lut_r_cen Ur8_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[0],sym_res_34_n[0],sym_res_33_n[0],sym_res_32_n[0] } ), .data_out( lut_val_8_n_0_pp[11:0]) ) ;
 defparam Ur8_n_0_pp.DATA_WIDTH = 12;
defparam Ur8_n_0_pp.C0 = 12'd                   0;
defparam Ur8_n_0_pp.C1 = 12'd                 154;
defparam Ur8_n_0_pp.C2 = 12'd                 377;
defparam Ur8_n_0_pp.C3 = 12'd                 531;
defparam Ur8_n_0_pp.C4 = 12'd                3846;
defparam Ur8_n_0_pp.C5 = 12'd                4000;
defparam Ur8_n_0_pp.C6 = 12'd                 127;
defparam Ur8_n_0_pp.C7 = 12'd                 281;
defparam Ur8_n_0_pp.C8 = 12'd                2476;
defparam Ur8_n_0_pp.C9 = 12'd                2630;
defparam Ur8_n_0_pp.CA = 12'd                2853;
defparam Ur8_n_0_pp.CB = 12'd                3007;
defparam Ur8_n_0_pp.CC = 12'd                2226;
defparam Ur8_n_0_pp.CD = 12'd                2380;
defparam Ur8_n_0_pp.CE = 12'd                2603;
defparam Ur8_n_0_pp.CF = 12'd                2757;
assign lut_val_8_n_0_pp[13] = lut_val_8_n_0_pp[11];
assign lut_val_8_n_0_pp[12] = lut_val_8_n_0_pp[11];
wire [13:0] lut_val_8_n_1_pp;
rom_lut_r_cen Ur8_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[1],sym_res_34_n[1],sym_res_33_n[1],sym_res_32_n[1] } ), .data_out( lut_val_8_n_1_pp[11:0]) ) ;
 defparam Ur8_n_1_pp.DATA_WIDTH = 12;
defparam Ur8_n_1_pp.C0 = 12'd                   0;
defparam Ur8_n_1_pp.C1 = 12'd                 154;
defparam Ur8_n_1_pp.C2 = 12'd                 377;
defparam Ur8_n_1_pp.C3 = 12'd                 531;
defparam Ur8_n_1_pp.C4 = 12'd                3846;
defparam Ur8_n_1_pp.C5 = 12'd                4000;
defparam Ur8_n_1_pp.C6 = 12'd                 127;
defparam Ur8_n_1_pp.C7 = 12'd                 281;
defparam Ur8_n_1_pp.C8 = 12'd                2476;
defparam Ur8_n_1_pp.C9 = 12'd                2630;
defparam Ur8_n_1_pp.CA = 12'd                2853;
defparam Ur8_n_1_pp.CB = 12'd                3007;
defparam Ur8_n_1_pp.CC = 12'd                2226;
defparam Ur8_n_1_pp.CD = 12'd                2380;
defparam Ur8_n_1_pp.CE = 12'd                2603;
defparam Ur8_n_1_pp.CF = 12'd                2757;
assign lut_val_8_n_1_pp[13] = lut_val_8_n_1_pp[11];
assign lut_val_8_n_1_pp[12] = lut_val_8_n_1_pp[11];
wire [13:0] lut_val_8_n_2_pp;
rom_lut_r_cen Ur8_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[2],sym_res_34_n[2],sym_res_33_n[2],sym_res_32_n[2] } ), .data_out( lut_val_8_n_2_pp[11:0]) ) ;
 defparam Ur8_n_2_pp.DATA_WIDTH = 12;
defparam Ur8_n_2_pp.C0 = 12'd                   0;
defparam Ur8_n_2_pp.C1 = 12'd                 154;
defparam Ur8_n_2_pp.C2 = 12'd                 377;
defparam Ur8_n_2_pp.C3 = 12'd                 531;
defparam Ur8_n_2_pp.C4 = 12'd                3846;
defparam Ur8_n_2_pp.C5 = 12'd                4000;
defparam Ur8_n_2_pp.C6 = 12'd                 127;
defparam Ur8_n_2_pp.C7 = 12'd                 281;
defparam Ur8_n_2_pp.C8 = 12'd                2476;
defparam Ur8_n_2_pp.C9 = 12'd                2630;
defparam Ur8_n_2_pp.CA = 12'd                2853;
defparam Ur8_n_2_pp.CB = 12'd                3007;
defparam Ur8_n_2_pp.CC = 12'd                2226;
defparam Ur8_n_2_pp.CD = 12'd                2380;
defparam Ur8_n_2_pp.CE = 12'd                2603;
defparam Ur8_n_2_pp.CF = 12'd                2757;
assign lut_val_8_n_2_pp[13] = lut_val_8_n_2_pp[11];
assign lut_val_8_n_2_pp[12] = lut_val_8_n_2_pp[11];
wire [13:0] lut_val_8_n_3_pp;
rom_lut_r_cen Ur8_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[3],sym_res_34_n[3],sym_res_33_n[3],sym_res_32_n[3] } ), .data_out( lut_val_8_n_3_pp[11:0]) ) ;
 defparam Ur8_n_3_pp.DATA_WIDTH = 12;
defparam Ur8_n_3_pp.C0 = 12'd                   0;
defparam Ur8_n_3_pp.C1 = 12'd                 154;
defparam Ur8_n_3_pp.C2 = 12'd                 377;
defparam Ur8_n_3_pp.C3 = 12'd                 531;
defparam Ur8_n_3_pp.C4 = 12'd                3846;
defparam Ur8_n_3_pp.C5 = 12'd                4000;
defparam Ur8_n_3_pp.C6 = 12'd                 127;
defparam Ur8_n_3_pp.C7 = 12'd                 281;
defparam Ur8_n_3_pp.C8 = 12'd                2476;
defparam Ur8_n_3_pp.C9 = 12'd                2630;
defparam Ur8_n_3_pp.CA = 12'd                2853;
defparam Ur8_n_3_pp.CB = 12'd                3007;
defparam Ur8_n_3_pp.CC = 12'd                2226;
defparam Ur8_n_3_pp.CD = 12'd                2380;
defparam Ur8_n_3_pp.CE = 12'd                2603;
defparam Ur8_n_3_pp.CF = 12'd                2757;
assign lut_val_8_n_3_pp[13] = lut_val_8_n_3_pp[11];
assign lut_val_8_n_3_pp[12] = lut_val_8_n_3_pp[11];
wire [13:0] lut_val_8_n_4_pp;
rom_lut_r_cen Ur8_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[4],sym_res_34_n[4],sym_res_33_n[4],sym_res_32_n[4] } ), .data_out( lut_val_8_n_4_pp[11:0]) ) ;
 defparam Ur8_n_4_pp.DATA_WIDTH = 12;
defparam Ur8_n_4_pp.C0 = 12'd                   0;
defparam Ur8_n_4_pp.C1 = 12'd                 154;
defparam Ur8_n_4_pp.C2 = 12'd                 377;
defparam Ur8_n_4_pp.C3 = 12'd                 531;
defparam Ur8_n_4_pp.C4 = 12'd                3846;
defparam Ur8_n_4_pp.C5 = 12'd                4000;
defparam Ur8_n_4_pp.C6 = 12'd                 127;
defparam Ur8_n_4_pp.C7 = 12'd                 281;
defparam Ur8_n_4_pp.C8 = 12'd                2476;
defparam Ur8_n_4_pp.C9 = 12'd                2630;
defparam Ur8_n_4_pp.CA = 12'd                2853;
defparam Ur8_n_4_pp.CB = 12'd                3007;
defparam Ur8_n_4_pp.CC = 12'd                2226;
defparam Ur8_n_4_pp.CD = 12'd                2380;
defparam Ur8_n_4_pp.CE = 12'd                2603;
defparam Ur8_n_4_pp.CF = 12'd                2757;
assign lut_val_8_n_4_pp[13] = lut_val_8_n_4_pp[11];
assign lut_val_8_n_4_pp[12] = lut_val_8_n_4_pp[11];
wire [13:0] lut_val_8_n_5_pp;
rom_lut_r_cen Ur8_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[5],sym_res_34_n[5],sym_res_33_n[5],sym_res_32_n[5] } ), .data_out( lut_val_8_n_5_pp[11:0]) ) ;
 defparam Ur8_n_5_pp.DATA_WIDTH = 12;
defparam Ur8_n_5_pp.C0 = 12'd                   0;
defparam Ur8_n_5_pp.C1 = 12'd                 154;
defparam Ur8_n_5_pp.C2 = 12'd                 377;
defparam Ur8_n_5_pp.C3 = 12'd                 531;
defparam Ur8_n_5_pp.C4 = 12'd                3846;
defparam Ur8_n_5_pp.C5 = 12'd                4000;
defparam Ur8_n_5_pp.C6 = 12'd                 127;
defparam Ur8_n_5_pp.C7 = 12'd                 281;
defparam Ur8_n_5_pp.C8 = 12'd                2476;
defparam Ur8_n_5_pp.C9 = 12'd                2630;
defparam Ur8_n_5_pp.CA = 12'd                2853;
defparam Ur8_n_5_pp.CB = 12'd                3007;
defparam Ur8_n_5_pp.CC = 12'd                2226;
defparam Ur8_n_5_pp.CD = 12'd                2380;
defparam Ur8_n_5_pp.CE = 12'd                2603;
defparam Ur8_n_5_pp.CF = 12'd                2757;
assign lut_val_8_n_5_pp[13] = lut_val_8_n_5_pp[11];
assign lut_val_8_n_5_pp[12] = lut_val_8_n_5_pp[11];
wire [13:0] lut_val_8_n_6_pp;
rom_lut_r_cen Ur8_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[6],sym_res_34_n[6],sym_res_33_n[6],sym_res_32_n[6] } ), .data_out( lut_val_8_n_6_pp[11:0]) ) ;
 defparam Ur8_n_6_pp.DATA_WIDTH = 12;
defparam Ur8_n_6_pp.C0 = 12'd                   0;
defparam Ur8_n_6_pp.C1 = 12'd                 154;
defparam Ur8_n_6_pp.C2 = 12'd                 377;
defparam Ur8_n_6_pp.C3 = 12'd                 531;
defparam Ur8_n_6_pp.C4 = 12'd                3846;
defparam Ur8_n_6_pp.C5 = 12'd                4000;
defparam Ur8_n_6_pp.C6 = 12'd                 127;
defparam Ur8_n_6_pp.C7 = 12'd                 281;
defparam Ur8_n_6_pp.C8 = 12'd                2476;
defparam Ur8_n_6_pp.C9 = 12'd                2630;
defparam Ur8_n_6_pp.CA = 12'd                2853;
defparam Ur8_n_6_pp.CB = 12'd                3007;
defparam Ur8_n_6_pp.CC = 12'd                2226;
defparam Ur8_n_6_pp.CD = 12'd                2380;
defparam Ur8_n_6_pp.CE = 12'd                2603;
defparam Ur8_n_6_pp.CF = 12'd                2757;
assign lut_val_8_n_6_pp[13] = lut_val_8_n_6_pp[11];
assign lut_val_8_n_6_pp[12] = lut_val_8_n_6_pp[11];
wire [13:0] lut_val_8_n_7_pp;
rom_lut_r_cen Ur8_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[7],sym_res_34_n[7],sym_res_33_n[7],sym_res_32_n[7] } ), .data_out( lut_val_8_n_7_pp[11:0]) ) ;
 defparam Ur8_n_7_pp.DATA_WIDTH = 12;
defparam Ur8_n_7_pp.C0 = 12'd                   0;
defparam Ur8_n_7_pp.C1 = 12'd                 154;
defparam Ur8_n_7_pp.C2 = 12'd                 377;
defparam Ur8_n_7_pp.C3 = 12'd                 531;
defparam Ur8_n_7_pp.C4 = 12'd                3846;
defparam Ur8_n_7_pp.C5 = 12'd                4000;
defparam Ur8_n_7_pp.C6 = 12'd                 127;
defparam Ur8_n_7_pp.C7 = 12'd                 281;
defparam Ur8_n_7_pp.C8 = 12'd                2476;
defparam Ur8_n_7_pp.C9 = 12'd                2630;
defparam Ur8_n_7_pp.CA = 12'd                2853;
defparam Ur8_n_7_pp.CB = 12'd                3007;
defparam Ur8_n_7_pp.CC = 12'd                2226;
defparam Ur8_n_7_pp.CD = 12'd                2380;
defparam Ur8_n_7_pp.CE = 12'd                2603;
defparam Ur8_n_7_pp.CF = 12'd                2757;
assign lut_val_8_n_7_pp[13] = lut_val_8_n_7_pp[11];
assign lut_val_8_n_7_pp[12] = lut_val_8_n_7_pp[11];
wire [13:0] lut_val_8_n_8_pp;
rom_lut_r_cen Ur8_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[8],sym_res_34_n[8],sym_res_33_n[8],sym_res_32_n[8] } ), .data_out( lut_val_8_n_8_pp[11:0]) ) ;
 defparam Ur8_n_8_pp.DATA_WIDTH = 12;
defparam Ur8_n_8_pp.C0 = 12'd                   0;
defparam Ur8_n_8_pp.C1 = 12'd                 154;
defparam Ur8_n_8_pp.C2 = 12'd                 377;
defparam Ur8_n_8_pp.C3 = 12'd                 531;
defparam Ur8_n_8_pp.C4 = 12'd                3846;
defparam Ur8_n_8_pp.C5 = 12'd                4000;
defparam Ur8_n_8_pp.C6 = 12'd                 127;
defparam Ur8_n_8_pp.C7 = 12'd                 281;
defparam Ur8_n_8_pp.C8 = 12'd                2476;
defparam Ur8_n_8_pp.C9 = 12'd                2630;
defparam Ur8_n_8_pp.CA = 12'd                2853;
defparam Ur8_n_8_pp.CB = 12'd                3007;
defparam Ur8_n_8_pp.CC = 12'd                2226;
defparam Ur8_n_8_pp.CD = 12'd                2380;
defparam Ur8_n_8_pp.CE = 12'd                2603;
defparam Ur8_n_8_pp.CF = 12'd                2757;
assign lut_val_8_n_8_pp[13] = lut_val_8_n_8_pp[11];
assign lut_val_8_n_8_pp[12] = lut_val_8_n_8_pp[11];
wire [13:0] lut_val_8_n_9_pp;
rom_lut_r_cen Ur8_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[9],sym_res_34_n[9],sym_res_33_n[9],sym_res_32_n[9] } ), .data_out( lut_val_8_n_9_pp[11:0]) ) ;
 defparam Ur8_n_9_pp.DATA_WIDTH = 12;
defparam Ur8_n_9_pp.C0 = 12'd                   0;
defparam Ur8_n_9_pp.C1 = 12'd                 154;
defparam Ur8_n_9_pp.C2 = 12'd                 377;
defparam Ur8_n_9_pp.C3 = 12'd                 531;
defparam Ur8_n_9_pp.C4 = 12'd                3846;
defparam Ur8_n_9_pp.C5 = 12'd                4000;
defparam Ur8_n_9_pp.C6 = 12'd                 127;
defparam Ur8_n_9_pp.C7 = 12'd                 281;
defparam Ur8_n_9_pp.C8 = 12'd                2476;
defparam Ur8_n_9_pp.C9 = 12'd                2630;
defparam Ur8_n_9_pp.CA = 12'd                2853;
defparam Ur8_n_9_pp.CB = 12'd                3007;
defparam Ur8_n_9_pp.CC = 12'd                2226;
defparam Ur8_n_9_pp.CD = 12'd                2380;
defparam Ur8_n_9_pp.CE = 12'd                2603;
defparam Ur8_n_9_pp.CF = 12'd                2757;
assign lut_val_8_n_9_pp[13] = lut_val_8_n_9_pp[11];
assign lut_val_8_n_9_pp[12] = lut_val_8_n_9_pp[11];
wire [13:0] lut_val_8_n_10_pp;
rom_lut_r_cen Ur8_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[10],sym_res_34_n[10],sym_res_33_n[10],sym_res_32_n[10] } ), .data_out( lut_val_8_n_10_pp[11:0]) ) ;
 defparam Ur8_n_10_pp.DATA_WIDTH = 12;
defparam Ur8_n_10_pp.C0 = 12'd                   0;
defparam Ur8_n_10_pp.C1 = 12'd                 154;
defparam Ur8_n_10_pp.C2 = 12'd                 377;
defparam Ur8_n_10_pp.C3 = 12'd                 531;
defparam Ur8_n_10_pp.C4 = 12'd                3846;
defparam Ur8_n_10_pp.C5 = 12'd                4000;
defparam Ur8_n_10_pp.C6 = 12'd                 127;
defparam Ur8_n_10_pp.C7 = 12'd                 281;
defparam Ur8_n_10_pp.C8 = 12'd                2476;
defparam Ur8_n_10_pp.C9 = 12'd                2630;
defparam Ur8_n_10_pp.CA = 12'd                2853;
defparam Ur8_n_10_pp.CB = 12'd                3007;
defparam Ur8_n_10_pp.CC = 12'd                2226;
defparam Ur8_n_10_pp.CD = 12'd                2380;
defparam Ur8_n_10_pp.CE = 12'd                2603;
defparam Ur8_n_10_pp.CF = 12'd                2757;
assign lut_val_8_n_10_pp[13] = lut_val_8_n_10_pp[11];
assign lut_val_8_n_10_pp[12] = lut_val_8_n_10_pp[11];
wire [13:0] lut_val_8_n_11_pp;
rom_lut_r_cen Ur8_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[11],sym_res_34_n[11],sym_res_33_n[11],sym_res_32_n[11] } ), .data_out( lut_val_8_n_11_pp[11:0]) ) ;
 defparam Ur8_n_11_pp.DATA_WIDTH = 12;
defparam Ur8_n_11_pp.C0 = 12'd                   0;
defparam Ur8_n_11_pp.C1 = 12'd                 154;
defparam Ur8_n_11_pp.C2 = 12'd                 377;
defparam Ur8_n_11_pp.C3 = 12'd                 531;
defparam Ur8_n_11_pp.C4 = 12'd                3846;
defparam Ur8_n_11_pp.C5 = 12'd                4000;
defparam Ur8_n_11_pp.C6 = 12'd                 127;
defparam Ur8_n_11_pp.C7 = 12'd                 281;
defparam Ur8_n_11_pp.C8 = 12'd                2476;
defparam Ur8_n_11_pp.C9 = 12'd                2630;
defparam Ur8_n_11_pp.CA = 12'd                2853;
defparam Ur8_n_11_pp.CB = 12'd                3007;
defparam Ur8_n_11_pp.CC = 12'd                2226;
defparam Ur8_n_11_pp.CD = 12'd                2380;
defparam Ur8_n_11_pp.CE = 12'd                2603;
defparam Ur8_n_11_pp.CF = 12'd                2757;
assign lut_val_8_n_11_pp[13] = lut_val_8_n_11_pp[11];
assign lut_val_8_n_11_pp[12] = lut_val_8_n_11_pp[11];
wire [13:0] lut_val_8_n_12_pp;
rom_lut_r_cen Ur8_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[12],sym_res_34_n[12],sym_res_33_n[12],sym_res_32_n[12] } ), .data_out( lut_val_8_n_12_pp[11:0]) ) ;
 defparam Ur8_n_12_pp.DATA_WIDTH = 12;
defparam Ur8_n_12_pp.C0 = 12'd                   0;
defparam Ur8_n_12_pp.C1 = 12'd                 154;
defparam Ur8_n_12_pp.C2 = 12'd                 377;
defparam Ur8_n_12_pp.C3 = 12'd                 531;
defparam Ur8_n_12_pp.C4 = 12'd                3846;
defparam Ur8_n_12_pp.C5 = 12'd                4000;
defparam Ur8_n_12_pp.C6 = 12'd                 127;
defparam Ur8_n_12_pp.C7 = 12'd                 281;
defparam Ur8_n_12_pp.C8 = 12'd                2476;
defparam Ur8_n_12_pp.C9 = 12'd                2630;
defparam Ur8_n_12_pp.CA = 12'd                2853;
defparam Ur8_n_12_pp.CB = 12'd                3007;
defparam Ur8_n_12_pp.CC = 12'd                2226;
defparam Ur8_n_12_pp.CD = 12'd                2380;
defparam Ur8_n_12_pp.CE = 12'd                2603;
defparam Ur8_n_12_pp.CF = 12'd                2757;
assign lut_val_8_n_12_pp[13] = lut_val_8_n_12_pp[11];
assign lut_val_8_n_12_pp[12] = lut_val_8_n_12_pp[11];
wire [13:0] lut_val_8_n_13_pp;
rom_lut_r_cen Ur8_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[13],sym_res_34_n[13],sym_res_33_n[13],sym_res_32_n[13] } ), .data_out( lut_val_8_n_13_pp[11:0]) ) ;
 defparam Ur8_n_13_pp.DATA_WIDTH = 12;
defparam Ur8_n_13_pp.C0 = 12'd                   0;
defparam Ur8_n_13_pp.C1 = 12'd                 154;
defparam Ur8_n_13_pp.C2 = 12'd                 377;
defparam Ur8_n_13_pp.C3 = 12'd                 531;
defparam Ur8_n_13_pp.C4 = 12'd                3846;
defparam Ur8_n_13_pp.C5 = 12'd                4000;
defparam Ur8_n_13_pp.C6 = 12'd                 127;
defparam Ur8_n_13_pp.C7 = 12'd                 281;
defparam Ur8_n_13_pp.C8 = 12'd                2476;
defparam Ur8_n_13_pp.C9 = 12'd                2630;
defparam Ur8_n_13_pp.CA = 12'd                2853;
defparam Ur8_n_13_pp.CB = 12'd                3007;
defparam Ur8_n_13_pp.CC = 12'd                2226;
defparam Ur8_n_13_pp.CD = 12'd                2380;
defparam Ur8_n_13_pp.CE = 12'd                2603;
defparam Ur8_n_13_pp.CF = 12'd                2757;
assign lut_val_8_n_13_pp[13] = lut_val_8_n_13_pp[11];
assign lut_val_8_n_13_pp[12] = lut_val_8_n_13_pp[11];
wire [13:0] lut_val_8_n_14_pp;
rom_lut_r_cen Ur8_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[14],sym_res_34_n[14],sym_res_33_n[14],sym_res_32_n[14] } ), .data_out( lut_val_8_n_14_pp[11:0]) ) ;
 defparam Ur8_n_14_pp.DATA_WIDTH = 12;
defparam Ur8_n_14_pp.C0 = 12'd                   0;
defparam Ur8_n_14_pp.C1 = 12'd                 154;
defparam Ur8_n_14_pp.C2 = 12'd                 377;
defparam Ur8_n_14_pp.C3 = 12'd                 531;
defparam Ur8_n_14_pp.C4 = 12'd                3846;
defparam Ur8_n_14_pp.C5 = 12'd                4000;
defparam Ur8_n_14_pp.C6 = 12'd                 127;
defparam Ur8_n_14_pp.C7 = 12'd                 281;
defparam Ur8_n_14_pp.C8 = 12'd                2476;
defparam Ur8_n_14_pp.C9 = 12'd                2630;
defparam Ur8_n_14_pp.CA = 12'd                2853;
defparam Ur8_n_14_pp.CB = 12'd                3007;
defparam Ur8_n_14_pp.CC = 12'd                2226;
defparam Ur8_n_14_pp.CD = 12'd                2380;
defparam Ur8_n_14_pp.CE = 12'd                2603;
defparam Ur8_n_14_pp.CF = 12'd                2757;
assign lut_val_8_n_14_pp[13] = lut_val_8_n_14_pp[11];
assign lut_val_8_n_14_pp[12] = lut_val_8_n_14_pp[11];
wire [13:0] lut_val_8_n_15_pp;
rom_lut_r_cen Ur8_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_35_n[15],sym_res_34_n[15],sym_res_33_n[15],sym_res_32_n[15] } ), .data_out( lut_val_8_n_15_pp[11:0]) ) ;
 defparam Ur8_n_15_pp.DATA_WIDTH = 12;
defparam Ur8_n_15_pp.C0 = 12'd                   0;
defparam Ur8_n_15_pp.C1 = 12'd                 154;
defparam Ur8_n_15_pp.C2 = 12'd                 377;
defparam Ur8_n_15_pp.C3 = 12'd                 531;
defparam Ur8_n_15_pp.C4 = 12'd                3846;
defparam Ur8_n_15_pp.C5 = 12'd                4000;
defparam Ur8_n_15_pp.C6 = 12'd                 127;
defparam Ur8_n_15_pp.C7 = 12'd                 281;
defparam Ur8_n_15_pp.C8 = 12'd                2476;
defparam Ur8_n_15_pp.C9 = 12'd                2630;
defparam Ur8_n_15_pp.CA = 12'd                2853;
defparam Ur8_n_15_pp.CB = 12'd                3007;
defparam Ur8_n_15_pp.CC = 12'd                2226;
defparam Ur8_n_15_pp.CD = 12'd                2380;
defparam Ur8_n_15_pp.CE = 12'd                2603;
defparam Ur8_n_15_pp.CF = 12'd                2757;
assign lut_val_8_n_15_pp[13] = lut_val_8_n_15_pp[11];
assign lut_val_8_n_15_pp[12] = lut_val_8_n_15_pp[11];
wire [13:0] lut_val_9_n_0_pp;
rom_lut_r_cen Ur9_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[0],sym_res_38_n[0],sym_res_37_n[0],sym_res_36_n[0] } ), .data_out( lut_val_9_n_0_pp[13:0]) ) ;
 defparam Ur9_n_0_pp.DATA_WIDTH = 14;
defparam Ur9_n_0_pp.C0 = 14'd                   0;
defparam Ur9_n_0_pp.C1 = 14'd               13749;
defparam Ur9_n_0_pp.C2 = 14'd               14320;
defparam Ur9_n_0_pp.C3 = 14'd               11685;
defparam Ur9_n_0_pp.C4 = 14'd                 232;
defparam Ur9_n_0_pp.C5 = 14'd               13981;
defparam Ur9_n_0_pp.C6 = 14'd               14552;
defparam Ur9_n_0_pp.C7 = 14'd               11917;
defparam Ur9_n_0_pp.C8 = 14'd                2911;
defparam Ur9_n_0_pp.C9 = 14'd                 276;
defparam Ur9_n_0_pp.CA = 14'd                 847;
defparam Ur9_n_0_pp.CB = 14'd               14596;
defparam Ur9_n_0_pp.CC = 14'd                3143;
defparam Ur9_n_0_pp.CD = 14'd                 508;
defparam Ur9_n_0_pp.CE = 14'd                1079;
defparam Ur9_n_0_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_1_pp;
rom_lut_r_cen Ur9_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[1],sym_res_38_n[1],sym_res_37_n[1],sym_res_36_n[1] } ), .data_out( lut_val_9_n_1_pp[13:0]) ) ;
 defparam Ur9_n_1_pp.DATA_WIDTH = 14;
defparam Ur9_n_1_pp.C0 = 14'd                   0;
defparam Ur9_n_1_pp.C1 = 14'd               13749;
defparam Ur9_n_1_pp.C2 = 14'd               14320;
defparam Ur9_n_1_pp.C3 = 14'd               11685;
defparam Ur9_n_1_pp.C4 = 14'd                 232;
defparam Ur9_n_1_pp.C5 = 14'd               13981;
defparam Ur9_n_1_pp.C6 = 14'd               14552;
defparam Ur9_n_1_pp.C7 = 14'd               11917;
defparam Ur9_n_1_pp.C8 = 14'd                2911;
defparam Ur9_n_1_pp.C9 = 14'd                 276;
defparam Ur9_n_1_pp.CA = 14'd                 847;
defparam Ur9_n_1_pp.CB = 14'd               14596;
defparam Ur9_n_1_pp.CC = 14'd                3143;
defparam Ur9_n_1_pp.CD = 14'd                 508;
defparam Ur9_n_1_pp.CE = 14'd                1079;
defparam Ur9_n_1_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_2_pp;
rom_lut_r_cen Ur9_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[2],sym_res_38_n[2],sym_res_37_n[2],sym_res_36_n[2] } ), .data_out( lut_val_9_n_2_pp[13:0]) ) ;
 defparam Ur9_n_2_pp.DATA_WIDTH = 14;
defparam Ur9_n_2_pp.C0 = 14'd                   0;
defparam Ur9_n_2_pp.C1 = 14'd               13749;
defparam Ur9_n_2_pp.C2 = 14'd               14320;
defparam Ur9_n_2_pp.C3 = 14'd               11685;
defparam Ur9_n_2_pp.C4 = 14'd                 232;
defparam Ur9_n_2_pp.C5 = 14'd               13981;
defparam Ur9_n_2_pp.C6 = 14'd               14552;
defparam Ur9_n_2_pp.C7 = 14'd               11917;
defparam Ur9_n_2_pp.C8 = 14'd                2911;
defparam Ur9_n_2_pp.C9 = 14'd                 276;
defparam Ur9_n_2_pp.CA = 14'd                 847;
defparam Ur9_n_2_pp.CB = 14'd               14596;
defparam Ur9_n_2_pp.CC = 14'd                3143;
defparam Ur9_n_2_pp.CD = 14'd                 508;
defparam Ur9_n_2_pp.CE = 14'd                1079;
defparam Ur9_n_2_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_3_pp;
rom_lut_r_cen Ur9_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[3],sym_res_38_n[3],sym_res_37_n[3],sym_res_36_n[3] } ), .data_out( lut_val_9_n_3_pp[13:0]) ) ;
 defparam Ur9_n_3_pp.DATA_WIDTH = 14;
defparam Ur9_n_3_pp.C0 = 14'd                   0;
defparam Ur9_n_3_pp.C1 = 14'd               13749;
defparam Ur9_n_3_pp.C2 = 14'd               14320;
defparam Ur9_n_3_pp.C3 = 14'd               11685;
defparam Ur9_n_3_pp.C4 = 14'd                 232;
defparam Ur9_n_3_pp.C5 = 14'd               13981;
defparam Ur9_n_3_pp.C6 = 14'd               14552;
defparam Ur9_n_3_pp.C7 = 14'd               11917;
defparam Ur9_n_3_pp.C8 = 14'd                2911;
defparam Ur9_n_3_pp.C9 = 14'd                 276;
defparam Ur9_n_3_pp.CA = 14'd                 847;
defparam Ur9_n_3_pp.CB = 14'd               14596;
defparam Ur9_n_3_pp.CC = 14'd                3143;
defparam Ur9_n_3_pp.CD = 14'd                 508;
defparam Ur9_n_3_pp.CE = 14'd                1079;
defparam Ur9_n_3_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_4_pp;
rom_lut_r_cen Ur9_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[4],sym_res_38_n[4],sym_res_37_n[4],sym_res_36_n[4] } ), .data_out( lut_val_9_n_4_pp[13:0]) ) ;
 defparam Ur9_n_4_pp.DATA_WIDTH = 14;
defparam Ur9_n_4_pp.C0 = 14'd                   0;
defparam Ur9_n_4_pp.C1 = 14'd               13749;
defparam Ur9_n_4_pp.C2 = 14'd               14320;
defparam Ur9_n_4_pp.C3 = 14'd               11685;
defparam Ur9_n_4_pp.C4 = 14'd                 232;
defparam Ur9_n_4_pp.C5 = 14'd               13981;
defparam Ur9_n_4_pp.C6 = 14'd               14552;
defparam Ur9_n_4_pp.C7 = 14'd               11917;
defparam Ur9_n_4_pp.C8 = 14'd                2911;
defparam Ur9_n_4_pp.C9 = 14'd                 276;
defparam Ur9_n_4_pp.CA = 14'd                 847;
defparam Ur9_n_4_pp.CB = 14'd               14596;
defparam Ur9_n_4_pp.CC = 14'd                3143;
defparam Ur9_n_4_pp.CD = 14'd                 508;
defparam Ur9_n_4_pp.CE = 14'd                1079;
defparam Ur9_n_4_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_5_pp;
rom_lut_r_cen Ur9_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[5],sym_res_38_n[5],sym_res_37_n[5],sym_res_36_n[5] } ), .data_out( lut_val_9_n_5_pp[13:0]) ) ;
 defparam Ur9_n_5_pp.DATA_WIDTH = 14;
defparam Ur9_n_5_pp.C0 = 14'd                   0;
defparam Ur9_n_5_pp.C1 = 14'd               13749;
defparam Ur9_n_5_pp.C2 = 14'd               14320;
defparam Ur9_n_5_pp.C3 = 14'd               11685;
defparam Ur9_n_5_pp.C4 = 14'd                 232;
defparam Ur9_n_5_pp.C5 = 14'd               13981;
defparam Ur9_n_5_pp.C6 = 14'd               14552;
defparam Ur9_n_5_pp.C7 = 14'd               11917;
defparam Ur9_n_5_pp.C8 = 14'd                2911;
defparam Ur9_n_5_pp.C9 = 14'd                 276;
defparam Ur9_n_5_pp.CA = 14'd                 847;
defparam Ur9_n_5_pp.CB = 14'd               14596;
defparam Ur9_n_5_pp.CC = 14'd                3143;
defparam Ur9_n_5_pp.CD = 14'd                 508;
defparam Ur9_n_5_pp.CE = 14'd                1079;
defparam Ur9_n_5_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_6_pp;
rom_lut_r_cen Ur9_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[6],sym_res_38_n[6],sym_res_37_n[6],sym_res_36_n[6] } ), .data_out( lut_val_9_n_6_pp[13:0]) ) ;
 defparam Ur9_n_6_pp.DATA_WIDTH = 14;
defparam Ur9_n_6_pp.C0 = 14'd                   0;
defparam Ur9_n_6_pp.C1 = 14'd               13749;
defparam Ur9_n_6_pp.C2 = 14'd               14320;
defparam Ur9_n_6_pp.C3 = 14'd               11685;
defparam Ur9_n_6_pp.C4 = 14'd                 232;
defparam Ur9_n_6_pp.C5 = 14'd               13981;
defparam Ur9_n_6_pp.C6 = 14'd               14552;
defparam Ur9_n_6_pp.C7 = 14'd               11917;
defparam Ur9_n_6_pp.C8 = 14'd                2911;
defparam Ur9_n_6_pp.C9 = 14'd                 276;
defparam Ur9_n_6_pp.CA = 14'd                 847;
defparam Ur9_n_6_pp.CB = 14'd               14596;
defparam Ur9_n_6_pp.CC = 14'd                3143;
defparam Ur9_n_6_pp.CD = 14'd                 508;
defparam Ur9_n_6_pp.CE = 14'd                1079;
defparam Ur9_n_6_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_7_pp;
rom_lut_r_cen Ur9_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[7],sym_res_38_n[7],sym_res_37_n[7],sym_res_36_n[7] } ), .data_out( lut_val_9_n_7_pp[13:0]) ) ;
 defparam Ur9_n_7_pp.DATA_WIDTH = 14;
defparam Ur9_n_7_pp.C0 = 14'd                   0;
defparam Ur9_n_7_pp.C1 = 14'd               13749;
defparam Ur9_n_7_pp.C2 = 14'd               14320;
defparam Ur9_n_7_pp.C3 = 14'd               11685;
defparam Ur9_n_7_pp.C4 = 14'd                 232;
defparam Ur9_n_7_pp.C5 = 14'd               13981;
defparam Ur9_n_7_pp.C6 = 14'd               14552;
defparam Ur9_n_7_pp.C7 = 14'd               11917;
defparam Ur9_n_7_pp.C8 = 14'd                2911;
defparam Ur9_n_7_pp.C9 = 14'd                 276;
defparam Ur9_n_7_pp.CA = 14'd                 847;
defparam Ur9_n_7_pp.CB = 14'd               14596;
defparam Ur9_n_7_pp.CC = 14'd                3143;
defparam Ur9_n_7_pp.CD = 14'd                 508;
defparam Ur9_n_7_pp.CE = 14'd                1079;
defparam Ur9_n_7_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_8_pp;
rom_lut_r_cen Ur9_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[8],sym_res_38_n[8],sym_res_37_n[8],sym_res_36_n[8] } ), .data_out( lut_val_9_n_8_pp[13:0]) ) ;
 defparam Ur9_n_8_pp.DATA_WIDTH = 14;
defparam Ur9_n_8_pp.C0 = 14'd                   0;
defparam Ur9_n_8_pp.C1 = 14'd               13749;
defparam Ur9_n_8_pp.C2 = 14'd               14320;
defparam Ur9_n_8_pp.C3 = 14'd               11685;
defparam Ur9_n_8_pp.C4 = 14'd                 232;
defparam Ur9_n_8_pp.C5 = 14'd               13981;
defparam Ur9_n_8_pp.C6 = 14'd               14552;
defparam Ur9_n_8_pp.C7 = 14'd               11917;
defparam Ur9_n_8_pp.C8 = 14'd                2911;
defparam Ur9_n_8_pp.C9 = 14'd                 276;
defparam Ur9_n_8_pp.CA = 14'd                 847;
defparam Ur9_n_8_pp.CB = 14'd               14596;
defparam Ur9_n_8_pp.CC = 14'd                3143;
defparam Ur9_n_8_pp.CD = 14'd                 508;
defparam Ur9_n_8_pp.CE = 14'd                1079;
defparam Ur9_n_8_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_9_pp;
rom_lut_r_cen Ur9_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[9],sym_res_38_n[9],sym_res_37_n[9],sym_res_36_n[9] } ), .data_out( lut_val_9_n_9_pp[13:0]) ) ;
 defparam Ur9_n_9_pp.DATA_WIDTH = 14;
defparam Ur9_n_9_pp.C0 = 14'd                   0;
defparam Ur9_n_9_pp.C1 = 14'd               13749;
defparam Ur9_n_9_pp.C2 = 14'd               14320;
defparam Ur9_n_9_pp.C3 = 14'd               11685;
defparam Ur9_n_9_pp.C4 = 14'd                 232;
defparam Ur9_n_9_pp.C5 = 14'd               13981;
defparam Ur9_n_9_pp.C6 = 14'd               14552;
defparam Ur9_n_9_pp.C7 = 14'd               11917;
defparam Ur9_n_9_pp.C8 = 14'd                2911;
defparam Ur9_n_9_pp.C9 = 14'd                 276;
defparam Ur9_n_9_pp.CA = 14'd                 847;
defparam Ur9_n_9_pp.CB = 14'd               14596;
defparam Ur9_n_9_pp.CC = 14'd                3143;
defparam Ur9_n_9_pp.CD = 14'd                 508;
defparam Ur9_n_9_pp.CE = 14'd                1079;
defparam Ur9_n_9_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_10_pp;
rom_lut_r_cen Ur9_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[10],sym_res_38_n[10],sym_res_37_n[10],sym_res_36_n[10] } ), .data_out( lut_val_9_n_10_pp[13:0]) ) ;
 defparam Ur9_n_10_pp.DATA_WIDTH = 14;
defparam Ur9_n_10_pp.C0 = 14'd                   0;
defparam Ur9_n_10_pp.C1 = 14'd               13749;
defparam Ur9_n_10_pp.C2 = 14'd               14320;
defparam Ur9_n_10_pp.C3 = 14'd               11685;
defparam Ur9_n_10_pp.C4 = 14'd                 232;
defparam Ur9_n_10_pp.C5 = 14'd               13981;
defparam Ur9_n_10_pp.C6 = 14'd               14552;
defparam Ur9_n_10_pp.C7 = 14'd               11917;
defparam Ur9_n_10_pp.C8 = 14'd                2911;
defparam Ur9_n_10_pp.C9 = 14'd                 276;
defparam Ur9_n_10_pp.CA = 14'd                 847;
defparam Ur9_n_10_pp.CB = 14'd               14596;
defparam Ur9_n_10_pp.CC = 14'd                3143;
defparam Ur9_n_10_pp.CD = 14'd                 508;
defparam Ur9_n_10_pp.CE = 14'd                1079;
defparam Ur9_n_10_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_11_pp;
rom_lut_r_cen Ur9_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[11],sym_res_38_n[11],sym_res_37_n[11],sym_res_36_n[11] } ), .data_out( lut_val_9_n_11_pp[13:0]) ) ;
 defparam Ur9_n_11_pp.DATA_WIDTH = 14;
defparam Ur9_n_11_pp.C0 = 14'd                   0;
defparam Ur9_n_11_pp.C1 = 14'd               13749;
defparam Ur9_n_11_pp.C2 = 14'd               14320;
defparam Ur9_n_11_pp.C3 = 14'd               11685;
defparam Ur9_n_11_pp.C4 = 14'd                 232;
defparam Ur9_n_11_pp.C5 = 14'd               13981;
defparam Ur9_n_11_pp.C6 = 14'd               14552;
defparam Ur9_n_11_pp.C7 = 14'd               11917;
defparam Ur9_n_11_pp.C8 = 14'd                2911;
defparam Ur9_n_11_pp.C9 = 14'd                 276;
defparam Ur9_n_11_pp.CA = 14'd                 847;
defparam Ur9_n_11_pp.CB = 14'd               14596;
defparam Ur9_n_11_pp.CC = 14'd                3143;
defparam Ur9_n_11_pp.CD = 14'd                 508;
defparam Ur9_n_11_pp.CE = 14'd                1079;
defparam Ur9_n_11_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_12_pp;
rom_lut_r_cen Ur9_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[12],sym_res_38_n[12],sym_res_37_n[12],sym_res_36_n[12] } ), .data_out( lut_val_9_n_12_pp[13:0]) ) ;
 defparam Ur9_n_12_pp.DATA_WIDTH = 14;
defparam Ur9_n_12_pp.C0 = 14'd                   0;
defparam Ur9_n_12_pp.C1 = 14'd               13749;
defparam Ur9_n_12_pp.C2 = 14'd               14320;
defparam Ur9_n_12_pp.C3 = 14'd               11685;
defparam Ur9_n_12_pp.C4 = 14'd                 232;
defparam Ur9_n_12_pp.C5 = 14'd               13981;
defparam Ur9_n_12_pp.C6 = 14'd               14552;
defparam Ur9_n_12_pp.C7 = 14'd               11917;
defparam Ur9_n_12_pp.C8 = 14'd                2911;
defparam Ur9_n_12_pp.C9 = 14'd                 276;
defparam Ur9_n_12_pp.CA = 14'd                 847;
defparam Ur9_n_12_pp.CB = 14'd               14596;
defparam Ur9_n_12_pp.CC = 14'd                3143;
defparam Ur9_n_12_pp.CD = 14'd                 508;
defparam Ur9_n_12_pp.CE = 14'd                1079;
defparam Ur9_n_12_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_13_pp;
rom_lut_r_cen Ur9_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[13],sym_res_38_n[13],sym_res_37_n[13],sym_res_36_n[13] } ), .data_out( lut_val_9_n_13_pp[13:0]) ) ;
 defparam Ur9_n_13_pp.DATA_WIDTH = 14;
defparam Ur9_n_13_pp.C0 = 14'd                   0;
defparam Ur9_n_13_pp.C1 = 14'd               13749;
defparam Ur9_n_13_pp.C2 = 14'd               14320;
defparam Ur9_n_13_pp.C3 = 14'd               11685;
defparam Ur9_n_13_pp.C4 = 14'd                 232;
defparam Ur9_n_13_pp.C5 = 14'd               13981;
defparam Ur9_n_13_pp.C6 = 14'd               14552;
defparam Ur9_n_13_pp.C7 = 14'd               11917;
defparam Ur9_n_13_pp.C8 = 14'd                2911;
defparam Ur9_n_13_pp.C9 = 14'd                 276;
defparam Ur9_n_13_pp.CA = 14'd                 847;
defparam Ur9_n_13_pp.CB = 14'd               14596;
defparam Ur9_n_13_pp.CC = 14'd                3143;
defparam Ur9_n_13_pp.CD = 14'd                 508;
defparam Ur9_n_13_pp.CE = 14'd                1079;
defparam Ur9_n_13_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_14_pp;
rom_lut_r_cen Ur9_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[14],sym_res_38_n[14],sym_res_37_n[14],sym_res_36_n[14] } ), .data_out( lut_val_9_n_14_pp[13:0]) ) ;
 defparam Ur9_n_14_pp.DATA_WIDTH = 14;
defparam Ur9_n_14_pp.C0 = 14'd                   0;
defparam Ur9_n_14_pp.C1 = 14'd               13749;
defparam Ur9_n_14_pp.C2 = 14'd               14320;
defparam Ur9_n_14_pp.C3 = 14'd               11685;
defparam Ur9_n_14_pp.C4 = 14'd                 232;
defparam Ur9_n_14_pp.C5 = 14'd               13981;
defparam Ur9_n_14_pp.C6 = 14'd               14552;
defparam Ur9_n_14_pp.C7 = 14'd               11917;
defparam Ur9_n_14_pp.C8 = 14'd                2911;
defparam Ur9_n_14_pp.C9 = 14'd                 276;
defparam Ur9_n_14_pp.CA = 14'd                 847;
defparam Ur9_n_14_pp.CB = 14'd               14596;
defparam Ur9_n_14_pp.CC = 14'd                3143;
defparam Ur9_n_14_pp.CD = 14'd                 508;
defparam Ur9_n_14_pp.CE = 14'd                1079;
defparam Ur9_n_14_pp.CF = 14'd               14828;
wire [13:0] lut_val_9_n_15_pp;
rom_lut_r_cen Ur9_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_39_n[15],sym_res_38_n[15],sym_res_37_n[15],sym_res_36_n[15] } ), .data_out( lut_val_9_n_15_pp[13:0]) ) ;
 defparam Ur9_n_15_pp.DATA_WIDTH = 14;
defparam Ur9_n_15_pp.C0 = 14'd                   0;
defparam Ur9_n_15_pp.C1 = 14'd               13749;
defparam Ur9_n_15_pp.C2 = 14'd               14320;
defparam Ur9_n_15_pp.C3 = 14'd               11685;
defparam Ur9_n_15_pp.C4 = 14'd                 232;
defparam Ur9_n_15_pp.C5 = 14'd               13981;
defparam Ur9_n_15_pp.C6 = 14'd               14552;
defparam Ur9_n_15_pp.C7 = 14'd               11917;
defparam Ur9_n_15_pp.C8 = 14'd                2911;
defparam Ur9_n_15_pp.C9 = 14'd                 276;
defparam Ur9_n_15_pp.CA = 14'd                 847;
defparam Ur9_n_15_pp.CB = 14'd               14596;
defparam Ur9_n_15_pp.CC = 14'd                3143;
defparam Ur9_n_15_pp.CD = 14'd                 508;
defparam Ur9_n_15_pp.CE = 14'd                1079;
defparam Ur9_n_15_pp.CF = 14'd               14828;
wire [13:0] lut_val_10_n_0_pp;
rom_lut_r_cen Ur10_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[0] } ), .data_out( lut_val_10_n_0_pp[12:0]) ) ;
 defparam Ur10_n_0_pp.DATA_WIDTH = 13;
defparam Ur10_n_0_pp.C0 = 13'd                   0;
defparam Ur10_n_0_pp.C1 = 13'd                4095;
defparam Ur10_n_0_pp.C2 = 13'd                   0;
defparam Ur10_n_0_pp.C3 = 13'd                4095;
defparam Ur10_n_0_pp.C4 = 13'd                   0;
defparam Ur10_n_0_pp.C5 = 13'd                4095;
defparam Ur10_n_0_pp.C6 = 13'd                   0;
defparam Ur10_n_0_pp.C7 = 13'd                4095;
defparam Ur10_n_0_pp.C8 = 13'd                   0;
defparam Ur10_n_0_pp.C9 = 13'd                4095;
defparam Ur10_n_0_pp.CA = 13'd                   0;
defparam Ur10_n_0_pp.CB = 13'd                4095;
defparam Ur10_n_0_pp.CC = 13'd                   0;
defparam Ur10_n_0_pp.CD = 13'd                4095;
defparam Ur10_n_0_pp.CE = 13'd                   0;
defparam Ur10_n_0_pp.CF = 13'd                4095;
assign lut_val_10_n_0_pp[13] = lut_val_10_n_0_pp[12];
wire [13:0] lut_val_10_n_1_pp;
rom_lut_r_cen Ur10_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[1] } ), .data_out( lut_val_10_n_1_pp[12:0]) ) ;
 defparam Ur10_n_1_pp.DATA_WIDTH = 13;
defparam Ur10_n_1_pp.C0 = 13'd                   0;
defparam Ur10_n_1_pp.C1 = 13'd                4095;
defparam Ur10_n_1_pp.C2 = 13'd                   0;
defparam Ur10_n_1_pp.C3 = 13'd                4095;
defparam Ur10_n_1_pp.C4 = 13'd                   0;
defparam Ur10_n_1_pp.C5 = 13'd                4095;
defparam Ur10_n_1_pp.C6 = 13'd                   0;
defparam Ur10_n_1_pp.C7 = 13'd                4095;
defparam Ur10_n_1_pp.C8 = 13'd                   0;
defparam Ur10_n_1_pp.C9 = 13'd                4095;
defparam Ur10_n_1_pp.CA = 13'd                   0;
defparam Ur10_n_1_pp.CB = 13'd                4095;
defparam Ur10_n_1_pp.CC = 13'd                   0;
defparam Ur10_n_1_pp.CD = 13'd                4095;
defparam Ur10_n_1_pp.CE = 13'd                   0;
defparam Ur10_n_1_pp.CF = 13'd                4095;
assign lut_val_10_n_1_pp[13] = lut_val_10_n_1_pp[12];
wire [13:0] lut_val_10_n_2_pp;
rom_lut_r_cen Ur10_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[2] } ), .data_out( lut_val_10_n_2_pp[12:0]) ) ;
 defparam Ur10_n_2_pp.DATA_WIDTH = 13;
defparam Ur10_n_2_pp.C0 = 13'd                   0;
defparam Ur10_n_2_pp.C1 = 13'd                4095;
defparam Ur10_n_2_pp.C2 = 13'd                   0;
defparam Ur10_n_2_pp.C3 = 13'd                4095;
defparam Ur10_n_2_pp.C4 = 13'd                   0;
defparam Ur10_n_2_pp.C5 = 13'd                4095;
defparam Ur10_n_2_pp.C6 = 13'd                   0;
defparam Ur10_n_2_pp.C7 = 13'd                4095;
defparam Ur10_n_2_pp.C8 = 13'd                   0;
defparam Ur10_n_2_pp.C9 = 13'd                4095;
defparam Ur10_n_2_pp.CA = 13'd                   0;
defparam Ur10_n_2_pp.CB = 13'd                4095;
defparam Ur10_n_2_pp.CC = 13'd                   0;
defparam Ur10_n_2_pp.CD = 13'd                4095;
defparam Ur10_n_2_pp.CE = 13'd                   0;
defparam Ur10_n_2_pp.CF = 13'd                4095;
assign lut_val_10_n_2_pp[13] = lut_val_10_n_2_pp[12];
wire [13:0] lut_val_10_n_3_pp;
rom_lut_r_cen Ur10_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[3] } ), .data_out( lut_val_10_n_3_pp[12:0]) ) ;
 defparam Ur10_n_3_pp.DATA_WIDTH = 13;
defparam Ur10_n_3_pp.C0 = 13'd                   0;
defparam Ur10_n_3_pp.C1 = 13'd                4095;
defparam Ur10_n_3_pp.C2 = 13'd                   0;
defparam Ur10_n_3_pp.C3 = 13'd                4095;
defparam Ur10_n_3_pp.C4 = 13'd                   0;
defparam Ur10_n_3_pp.C5 = 13'd                4095;
defparam Ur10_n_3_pp.C6 = 13'd                   0;
defparam Ur10_n_3_pp.C7 = 13'd                4095;
defparam Ur10_n_3_pp.C8 = 13'd                   0;
defparam Ur10_n_3_pp.C9 = 13'd                4095;
defparam Ur10_n_3_pp.CA = 13'd                   0;
defparam Ur10_n_3_pp.CB = 13'd                4095;
defparam Ur10_n_3_pp.CC = 13'd                   0;
defparam Ur10_n_3_pp.CD = 13'd                4095;
defparam Ur10_n_3_pp.CE = 13'd                   0;
defparam Ur10_n_3_pp.CF = 13'd                4095;
assign lut_val_10_n_3_pp[13] = lut_val_10_n_3_pp[12];
wire [13:0] lut_val_10_n_4_pp;
rom_lut_r_cen Ur10_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[4] } ), .data_out( lut_val_10_n_4_pp[12:0]) ) ;
 defparam Ur10_n_4_pp.DATA_WIDTH = 13;
defparam Ur10_n_4_pp.C0 = 13'd                   0;
defparam Ur10_n_4_pp.C1 = 13'd                4095;
defparam Ur10_n_4_pp.C2 = 13'd                   0;
defparam Ur10_n_4_pp.C3 = 13'd                4095;
defparam Ur10_n_4_pp.C4 = 13'd                   0;
defparam Ur10_n_4_pp.C5 = 13'd                4095;
defparam Ur10_n_4_pp.C6 = 13'd                   0;
defparam Ur10_n_4_pp.C7 = 13'd                4095;
defparam Ur10_n_4_pp.C8 = 13'd                   0;
defparam Ur10_n_4_pp.C9 = 13'd                4095;
defparam Ur10_n_4_pp.CA = 13'd                   0;
defparam Ur10_n_4_pp.CB = 13'd                4095;
defparam Ur10_n_4_pp.CC = 13'd                   0;
defparam Ur10_n_4_pp.CD = 13'd                4095;
defparam Ur10_n_4_pp.CE = 13'd                   0;
defparam Ur10_n_4_pp.CF = 13'd                4095;
assign lut_val_10_n_4_pp[13] = lut_val_10_n_4_pp[12];
wire [13:0] lut_val_10_n_5_pp;
rom_lut_r_cen Ur10_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[5] } ), .data_out( lut_val_10_n_5_pp[12:0]) ) ;
 defparam Ur10_n_5_pp.DATA_WIDTH = 13;
defparam Ur10_n_5_pp.C0 = 13'd                   0;
defparam Ur10_n_5_pp.C1 = 13'd                4095;
defparam Ur10_n_5_pp.C2 = 13'd                   0;
defparam Ur10_n_5_pp.C3 = 13'd                4095;
defparam Ur10_n_5_pp.C4 = 13'd                   0;
defparam Ur10_n_5_pp.C5 = 13'd                4095;
defparam Ur10_n_5_pp.C6 = 13'd                   0;
defparam Ur10_n_5_pp.C7 = 13'd                4095;
defparam Ur10_n_5_pp.C8 = 13'd                   0;
defparam Ur10_n_5_pp.C9 = 13'd                4095;
defparam Ur10_n_5_pp.CA = 13'd                   0;
defparam Ur10_n_5_pp.CB = 13'd                4095;
defparam Ur10_n_5_pp.CC = 13'd                   0;
defparam Ur10_n_5_pp.CD = 13'd                4095;
defparam Ur10_n_5_pp.CE = 13'd                   0;
defparam Ur10_n_5_pp.CF = 13'd                4095;
assign lut_val_10_n_5_pp[13] = lut_val_10_n_5_pp[12];
wire [13:0] lut_val_10_n_6_pp;
rom_lut_r_cen Ur10_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[6] } ), .data_out( lut_val_10_n_6_pp[12:0]) ) ;
 defparam Ur10_n_6_pp.DATA_WIDTH = 13;
defparam Ur10_n_6_pp.C0 = 13'd                   0;
defparam Ur10_n_6_pp.C1 = 13'd                4095;
defparam Ur10_n_6_pp.C2 = 13'd                   0;
defparam Ur10_n_6_pp.C3 = 13'd                4095;
defparam Ur10_n_6_pp.C4 = 13'd                   0;
defparam Ur10_n_6_pp.C5 = 13'd                4095;
defparam Ur10_n_6_pp.C6 = 13'd                   0;
defparam Ur10_n_6_pp.C7 = 13'd                4095;
defparam Ur10_n_6_pp.C8 = 13'd                   0;
defparam Ur10_n_6_pp.C9 = 13'd                4095;
defparam Ur10_n_6_pp.CA = 13'd                   0;
defparam Ur10_n_6_pp.CB = 13'd                4095;
defparam Ur10_n_6_pp.CC = 13'd                   0;
defparam Ur10_n_6_pp.CD = 13'd                4095;
defparam Ur10_n_6_pp.CE = 13'd                   0;
defparam Ur10_n_6_pp.CF = 13'd                4095;
assign lut_val_10_n_6_pp[13] = lut_val_10_n_6_pp[12];
wire [13:0] lut_val_10_n_7_pp;
rom_lut_r_cen Ur10_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[7] } ), .data_out( lut_val_10_n_7_pp[12:0]) ) ;
 defparam Ur10_n_7_pp.DATA_WIDTH = 13;
defparam Ur10_n_7_pp.C0 = 13'd                   0;
defparam Ur10_n_7_pp.C1 = 13'd                4095;
defparam Ur10_n_7_pp.C2 = 13'd                   0;
defparam Ur10_n_7_pp.C3 = 13'd                4095;
defparam Ur10_n_7_pp.C4 = 13'd                   0;
defparam Ur10_n_7_pp.C5 = 13'd                4095;
defparam Ur10_n_7_pp.C6 = 13'd                   0;
defparam Ur10_n_7_pp.C7 = 13'd                4095;
defparam Ur10_n_7_pp.C8 = 13'd                   0;
defparam Ur10_n_7_pp.C9 = 13'd                4095;
defparam Ur10_n_7_pp.CA = 13'd                   0;
defparam Ur10_n_7_pp.CB = 13'd                4095;
defparam Ur10_n_7_pp.CC = 13'd                   0;
defparam Ur10_n_7_pp.CD = 13'd                4095;
defparam Ur10_n_7_pp.CE = 13'd                   0;
defparam Ur10_n_7_pp.CF = 13'd                4095;
assign lut_val_10_n_7_pp[13] = lut_val_10_n_7_pp[12];
wire [13:0] lut_val_10_n_8_pp;
rom_lut_r_cen Ur10_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[8] } ), .data_out( lut_val_10_n_8_pp[12:0]) ) ;
 defparam Ur10_n_8_pp.DATA_WIDTH = 13;
defparam Ur10_n_8_pp.C0 = 13'd                   0;
defparam Ur10_n_8_pp.C1 = 13'd                4095;
defparam Ur10_n_8_pp.C2 = 13'd                   0;
defparam Ur10_n_8_pp.C3 = 13'd                4095;
defparam Ur10_n_8_pp.C4 = 13'd                   0;
defparam Ur10_n_8_pp.C5 = 13'd                4095;
defparam Ur10_n_8_pp.C6 = 13'd                   0;
defparam Ur10_n_8_pp.C7 = 13'd                4095;
defparam Ur10_n_8_pp.C8 = 13'd                   0;
defparam Ur10_n_8_pp.C9 = 13'd                4095;
defparam Ur10_n_8_pp.CA = 13'd                   0;
defparam Ur10_n_8_pp.CB = 13'd                4095;
defparam Ur10_n_8_pp.CC = 13'd                   0;
defparam Ur10_n_8_pp.CD = 13'd                4095;
defparam Ur10_n_8_pp.CE = 13'd                   0;
defparam Ur10_n_8_pp.CF = 13'd                4095;
assign lut_val_10_n_8_pp[13] = lut_val_10_n_8_pp[12];
wire [13:0] lut_val_10_n_9_pp;
rom_lut_r_cen Ur10_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[9] } ), .data_out( lut_val_10_n_9_pp[12:0]) ) ;
 defparam Ur10_n_9_pp.DATA_WIDTH = 13;
defparam Ur10_n_9_pp.C0 = 13'd                   0;
defparam Ur10_n_9_pp.C1 = 13'd                4095;
defparam Ur10_n_9_pp.C2 = 13'd                   0;
defparam Ur10_n_9_pp.C3 = 13'd                4095;
defparam Ur10_n_9_pp.C4 = 13'd                   0;
defparam Ur10_n_9_pp.C5 = 13'd                4095;
defparam Ur10_n_9_pp.C6 = 13'd                   0;
defparam Ur10_n_9_pp.C7 = 13'd                4095;
defparam Ur10_n_9_pp.C8 = 13'd                   0;
defparam Ur10_n_9_pp.C9 = 13'd                4095;
defparam Ur10_n_9_pp.CA = 13'd                   0;
defparam Ur10_n_9_pp.CB = 13'd                4095;
defparam Ur10_n_9_pp.CC = 13'd                   0;
defparam Ur10_n_9_pp.CD = 13'd                4095;
defparam Ur10_n_9_pp.CE = 13'd                   0;
defparam Ur10_n_9_pp.CF = 13'd                4095;
assign lut_val_10_n_9_pp[13] = lut_val_10_n_9_pp[12];
wire [13:0] lut_val_10_n_10_pp;
rom_lut_r_cen Ur10_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[10] } ), .data_out( lut_val_10_n_10_pp[12:0]) ) ;
 defparam Ur10_n_10_pp.DATA_WIDTH = 13;
defparam Ur10_n_10_pp.C0 = 13'd                   0;
defparam Ur10_n_10_pp.C1 = 13'd                4095;
defparam Ur10_n_10_pp.C2 = 13'd                   0;
defparam Ur10_n_10_pp.C3 = 13'd                4095;
defparam Ur10_n_10_pp.C4 = 13'd                   0;
defparam Ur10_n_10_pp.C5 = 13'd                4095;
defparam Ur10_n_10_pp.C6 = 13'd                   0;
defparam Ur10_n_10_pp.C7 = 13'd                4095;
defparam Ur10_n_10_pp.C8 = 13'd                   0;
defparam Ur10_n_10_pp.C9 = 13'd                4095;
defparam Ur10_n_10_pp.CA = 13'd                   0;
defparam Ur10_n_10_pp.CB = 13'd                4095;
defparam Ur10_n_10_pp.CC = 13'd                   0;
defparam Ur10_n_10_pp.CD = 13'd                4095;
defparam Ur10_n_10_pp.CE = 13'd                   0;
defparam Ur10_n_10_pp.CF = 13'd                4095;
assign lut_val_10_n_10_pp[13] = lut_val_10_n_10_pp[12];
wire [13:0] lut_val_10_n_11_pp;
rom_lut_r_cen Ur10_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[11] } ), .data_out( lut_val_10_n_11_pp[12:0]) ) ;
 defparam Ur10_n_11_pp.DATA_WIDTH = 13;
defparam Ur10_n_11_pp.C0 = 13'd                   0;
defparam Ur10_n_11_pp.C1 = 13'd                4095;
defparam Ur10_n_11_pp.C2 = 13'd                   0;
defparam Ur10_n_11_pp.C3 = 13'd                4095;
defparam Ur10_n_11_pp.C4 = 13'd                   0;
defparam Ur10_n_11_pp.C5 = 13'd                4095;
defparam Ur10_n_11_pp.C6 = 13'd                   0;
defparam Ur10_n_11_pp.C7 = 13'd                4095;
defparam Ur10_n_11_pp.C8 = 13'd                   0;
defparam Ur10_n_11_pp.C9 = 13'd                4095;
defparam Ur10_n_11_pp.CA = 13'd                   0;
defparam Ur10_n_11_pp.CB = 13'd                4095;
defparam Ur10_n_11_pp.CC = 13'd                   0;
defparam Ur10_n_11_pp.CD = 13'd                4095;
defparam Ur10_n_11_pp.CE = 13'd                   0;
defparam Ur10_n_11_pp.CF = 13'd                4095;
assign lut_val_10_n_11_pp[13] = lut_val_10_n_11_pp[12];
wire [13:0] lut_val_10_n_12_pp;
rom_lut_r_cen Ur10_n_12_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[12] } ), .data_out( lut_val_10_n_12_pp[12:0]) ) ;
 defparam Ur10_n_12_pp.DATA_WIDTH = 13;
defparam Ur10_n_12_pp.C0 = 13'd                   0;
defparam Ur10_n_12_pp.C1 = 13'd                4095;
defparam Ur10_n_12_pp.C2 = 13'd                   0;
defparam Ur10_n_12_pp.C3 = 13'd                4095;
defparam Ur10_n_12_pp.C4 = 13'd                   0;
defparam Ur10_n_12_pp.C5 = 13'd                4095;
defparam Ur10_n_12_pp.C6 = 13'd                   0;
defparam Ur10_n_12_pp.C7 = 13'd                4095;
defparam Ur10_n_12_pp.C8 = 13'd                   0;
defparam Ur10_n_12_pp.C9 = 13'd                4095;
defparam Ur10_n_12_pp.CA = 13'd                   0;
defparam Ur10_n_12_pp.CB = 13'd                4095;
defparam Ur10_n_12_pp.CC = 13'd                   0;
defparam Ur10_n_12_pp.CD = 13'd                4095;
defparam Ur10_n_12_pp.CE = 13'd                   0;
defparam Ur10_n_12_pp.CF = 13'd                4095;
assign lut_val_10_n_12_pp[13] = lut_val_10_n_12_pp[12];
wire [13:0] lut_val_10_n_13_pp;
rom_lut_r_cen Ur10_n_13_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[13] } ), .data_out( lut_val_10_n_13_pp[12:0]) ) ;
 defparam Ur10_n_13_pp.DATA_WIDTH = 13;
defparam Ur10_n_13_pp.C0 = 13'd                   0;
defparam Ur10_n_13_pp.C1 = 13'd                4095;
defparam Ur10_n_13_pp.C2 = 13'd                   0;
defparam Ur10_n_13_pp.C3 = 13'd                4095;
defparam Ur10_n_13_pp.C4 = 13'd                   0;
defparam Ur10_n_13_pp.C5 = 13'd                4095;
defparam Ur10_n_13_pp.C6 = 13'd                   0;
defparam Ur10_n_13_pp.C7 = 13'd                4095;
defparam Ur10_n_13_pp.C8 = 13'd                   0;
defparam Ur10_n_13_pp.C9 = 13'd                4095;
defparam Ur10_n_13_pp.CA = 13'd                   0;
defparam Ur10_n_13_pp.CB = 13'd                4095;
defparam Ur10_n_13_pp.CC = 13'd                   0;
defparam Ur10_n_13_pp.CD = 13'd                4095;
defparam Ur10_n_13_pp.CE = 13'd                   0;
defparam Ur10_n_13_pp.CF = 13'd                4095;
assign lut_val_10_n_13_pp[13] = lut_val_10_n_13_pp[12];
wire [13:0] lut_val_10_n_14_pp;
rom_lut_r_cen Ur10_n_14_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[14] } ), .data_out( lut_val_10_n_14_pp[12:0]) ) ;
 defparam Ur10_n_14_pp.DATA_WIDTH = 13;
defparam Ur10_n_14_pp.C0 = 13'd                   0;
defparam Ur10_n_14_pp.C1 = 13'd                4095;
defparam Ur10_n_14_pp.C2 = 13'd                   0;
defparam Ur10_n_14_pp.C3 = 13'd                4095;
defparam Ur10_n_14_pp.C4 = 13'd                   0;
defparam Ur10_n_14_pp.C5 = 13'd                4095;
defparam Ur10_n_14_pp.C6 = 13'd                   0;
defparam Ur10_n_14_pp.C7 = 13'd                4095;
defparam Ur10_n_14_pp.C8 = 13'd                   0;
defparam Ur10_n_14_pp.C9 = 13'd                4095;
defparam Ur10_n_14_pp.CA = 13'd                   0;
defparam Ur10_n_14_pp.CB = 13'd                4095;
defparam Ur10_n_14_pp.CC = 13'd                   0;
defparam Ur10_n_14_pp.CD = 13'd                4095;
defparam Ur10_n_14_pp.CE = 13'd                   0;
defparam Ur10_n_14_pp.CF = 13'd                4095;
assign lut_val_10_n_14_pp[13] = lut_val_10_n_14_pp[12];
wire [13:0] lut_val_10_n_15_pp;
rom_lut_r_cen Ur10_n_15_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,addr_low,sym_res_40_n[15] } ), .data_out( lut_val_10_n_15_pp[12:0]) ) ;
 defparam Ur10_n_15_pp.DATA_WIDTH = 13;
defparam Ur10_n_15_pp.C0 = 13'd                   0;
defparam Ur10_n_15_pp.C1 = 13'd                4095;
defparam Ur10_n_15_pp.C2 = 13'd                   0;
defparam Ur10_n_15_pp.C3 = 13'd                4095;
defparam Ur10_n_15_pp.C4 = 13'd                   0;
defparam Ur10_n_15_pp.C5 = 13'd                4095;
defparam Ur10_n_15_pp.C6 = 13'd                   0;
defparam Ur10_n_15_pp.C7 = 13'd                4095;
defparam Ur10_n_15_pp.C8 = 13'd                   0;
defparam Ur10_n_15_pp.C9 = 13'd                4095;
defparam Ur10_n_15_pp.CA = 13'd                   0;
defparam Ur10_n_15_pp.CB = 13'd                4095;
defparam Ur10_n_15_pp.CC = 13'd                   0;
defparam Ur10_n_15_pp.CD = 13'd                4095;
defparam Ur10_n_15_pp.CE = 13'd                   0;
defparam Ur10_n_15_pp.CF = 13'd                4095;
assign lut_val_10_n_15_pp[13] = lut_val_10_n_15_pp[12];
wire [28:0] lut_0_bit_0_fill;
wire [28:0] lut_0_bit_1_fill;
wire [28:0] lut_0_bit_2_fill;
wire [28:0] lut_0_bit_3_fill;
wire [28:0] lut_0_bit_4_fill;
wire [28:0] lut_0_bit_5_fill;
wire [28:0] lut_0_bit_6_fill;
wire [28:0] lut_0_bit_7_fill;
wire [28:0] lut_0_bit_8_fill;
wire [28:0] lut_0_bit_9_fill;
wire [28:0] lut_0_bit_10_fill;
wire [28:0] lut_0_bit_11_fill;
wire [28:0] lut_0_bit_12_fill;
wire [28:0] lut_0_bit_13_fill;
wire [28:0] lut_0_bit_14_fill;
wire [28:0] lut_0_bit_15_fill;
assign lut_0_bit_0_fill = {lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13], lut_val_0_n_0_pp[13],  lut_val_0_n_0_pp };
assign lut_0_bit_1_fill = {lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13], lut_val_0_n_1_pp[13],  lut_val_0_n_1_pp, 1'd0 };
assign lut_0_bit_2_fill = {lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13], lut_val_0_n_2_pp[13],  lut_val_0_n_2_pp, 2'd0 };
assign lut_0_bit_3_fill = {lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13], lut_val_0_n_3_pp[13],  lut_val_0_n_3_pp, 3'd0 };
assign lut_0_bit_4_fill = {lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13], lut_val_0_n_4_pp[13],  lut_val_0_n_4_pp, 4'd0 };
assign lut_0_bit_5_fill = {lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13], lut_val_0_n_5_pp[13],  lut_val_0_n_5_pp, 5'd0 };
assign lut_0_bit_6_fill = {lut_val_0_n_6_pp[13], lut_val_0_n_6_pp[13], lut_val_0_n_6_pp[13], lut_val_0_n_6_pp[13], lut_val_0_n_6_pp[13], lut_val_0_n_6_pp[13], lut_val_0_n_6_pp[13], lut_val_0_n_6_pp[13], lut_val_0_n_6_pp[13],  lut_val_0_n_6_pp, 6'd0 };
assign lut_0_bit_7_fill = {lut_val_0_n_7_pp[13], lut_val_0_n_7_pp[13], lut_val_0_n_7_pp[13], lut_val_0_n_7_pp[13], lut_val_0_n_7_pp[13], lut_val_0_n_7_pp[13], lut_val_0_n_7_pp[13], lut_val_0_n_7_pp[13],  lut_val_0_n_7_pp, 7'd0 };
assign lut_0_bit_8_fill = {lut_val_0_n_8_pp[13], lut_val_0_n_8_pp[13], lut_val_0_n_8_pp[13], lut_val_0_n_8_pp[13], lut_val_0_n_8_pp[13], lut_val_0_n_8_pp[13], lut_val_0_n_8_pp[13],  lut_val_0_n_8_pp, 8'd0 };
assign lut_0_bit_9_fill = {lut_val_0_n_9_pp[13], lut_val_0_n_9_pp[13], lut_val_0_n_9_pp[13], lut_val_0_n_9_pp[13], lut_val_0_n_9_pp[13], lut_val_0_n_9_pp[13],  lut_val_0_n_9_pp, 9'd0 };
assign lut_0_bit_10_fill = {lut_val_0_n_10_pp[13], lut_val_0_n_10_pp[13], lut_val_0_n_10_pp[13], lut_val_0_n_10_pp[13], lut_val_0_n_10_pp[13],  lut_val_0_n_10_pp, 10'd0 };
assign lut_0_bit_11_fill = {lut_val_0_n_11_pp[13], lut_val_0_n_11_pp[13], lut_val_0_n_11_pp[13], lut_val_0_n_11_pp[13],  lut_val_0_n_11_pp, 11'd0 };
assign lut_0_bit_12_fill = {lut_val_0_n_12_pp[13], lut_val_0_n_12_pp[13], lut_val_0_n_12_pp[13],  lut_val_0_n_12_pp, 12'd0 };
assign lut_0_bit_13_fill = {lut_val_0_n_13_pp[13], lut_val_0_n_13_pp[13],  lut_val_0_n_13_pp, 13'd0 };
assign lut_0_bit_14_fill = {lut_val_0_n_14_pp[13],  lut_val_0_n_14_pp, 14'd0 };
assign lut_0_bit_15_fill = { lut_val_0_n_15_pp, 15'd0 };
wire [29:0] tree_0_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_0_fill), .bin(lut_0_bit_1_fill), .res(tree_0_pp_l_0_n_0_n) );
defparam Uadd_0_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_0_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_0_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_2_fill), .bin(lut_0_bit_3_fill), .res(tree_0_pp_l_0_n_1_n) );
defparam Uadd_0_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_0_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_0_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_4_fill), .bin(lut_0_bit_5_fill), .res(tree_0_pp_l_0_n_2_n) );
defparam Uadd_0_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_0_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_0_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_6_fill), .bin(lut_0_bit_7_fill), .res(tree_0_pp_l_0_n_3_n) );
defparam Uadd_0_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_0_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_0_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_8_fill), .bin(lut_0_bit_9_fill), .res(tree_0_pp_l_0_n_4_n) );
defparam Uadd_0_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_0_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_0_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_10_fill), .bin(lut_0_bit_11_fill), .res(tree_0_pp_l_0_n_5_n) );
defparam Uadd_0_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_0_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_0_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_12_fill), .bin(lut_0_bit_13_fill), .res(tree_0_pp_l_0_n_6_n) );
defparam Uadd_0_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_0_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_0_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_14_fill), .bin(lut_0_bit_15_fill), .res(tree_0_pp_l_0_n_7_n) );
defparam Uadd_0_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_0_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_0_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_0_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_0_n_0_n), .bin(tree_0_pp_l_0_n_1_n), .res(tree_0_pp_l_1_n_0_n) );
defparam Uadd_0_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_0_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_0_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_0_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_0_n_2_n), .bin(tree_0_pp_l_0_n_3_n), .res(tree_0_pp_l_1_n_1_n) );
defparam Uadd_0_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_0_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_0_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_0_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_0_n_4_n), .bin(tree_0_pp_l_0_n_5_n), .res(tree_0_pp_l_1_n_2_n) );
defparam Uadd_0_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_0_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_0_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_0_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_0_n_6_n), .bin(tree_0_pp_l_0_n_7_n), .res(tree_0_pp_l_1_n_3_n) );
defparam Uadd_0_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_0_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_0_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_0_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_1_n_0_n), .bin(tree_0_pp_l_1_n_1_n), .res(tree_0_pp_l_2_n_0_n) );
defparam Uadd_0_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_0_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_0_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_0_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_1_n_2_n), .bin(tree_0_pp_l_1_n_3_n), .res(tree_0_pp_l_2_n_1_n) );
defparam Uadd_0_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_0_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_0_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_0_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_2_n_0_n), .bin(tree_0_pp_l_2_n_1_n), .res(tree_0_pp_l_3_n_0_n) );
defparam Uadd_0_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_0_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_0_n;
assign lut_val_0_n=tree_0_pp_l_3_n_0_n;
wire [28:0] lut_1_bit_0_fill;
wire [28:0] lut_1_bit_1_fill;
wire [28:0] lut_1_bit_2_fill;
wire [28:0] lut_1_bit_3_fill;
wire [28:0] lut_1_bit_4_fill;
wire [28:0] lut_1_bit_5_fill;
wire [28:0] lut_1_bit_6_fill;
wire [28:0] lut_1_bit_7_fill;
wire [28:0] lut_1_bit_8_fill;
wire [28:0] lut_1_bit_9_fill;
wire [28:0] lut_1_bit_10_fill;
wire [28:0] lut_1_bit_11_fill;
wire [28:0] lut_1_bit_12_fill;
wire [28:0] lut_1_bit_13_fill;
wire [28:0] lut_1_bit_14_fill;
wire [28:0] lut_1_bit_15_fill;
assign lut_1_bit_0_fill = {lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13], lut_val_1_n_0_pp[13],  lut_val_1_n_0_pp };
assign lut_1_bit_1_fill = {lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13], lut_val_1_n_1_pp[13],  lut_val_1_n_1_pp, 1'd0 };
assign lut_1_bit_2_fill = {lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13], lut_val_1_n_2_pp[13],  lut_val_1_n_2_pp, 2'd0 };
assign lut_1_bit_3_fill = {lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13], lut_val_1_n_3_pp[13],  lut_val_1_n_3_pp, 3'd0 };
assign lut_1_bit_4_fill = {lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13], lut_val_1_n_4_pp[13],  lut_val_1_n_4_pp, 4'd0 };
assign lut_1_bit_5_fill = {lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13], lut_val_1_n_5_pp[13],  lut_val_1_n_5_pp, 5'd0 };
assign lut_1_bit_6_fill = {lut_val_1_n_6_pp[13], lut_val_1_n_6_pp[13], lut_val_1_n_6_pp[13], lut_val_1_n_6_pp[13], lut_val_1_n_6_pp[13], lut_val_1_n_6_pp[13], lut_val_1_n_6_pp[13], lut_val_1_n_6_pp[13], lut_val_1_n_6_pp[13],  lut_val_1_n_6_pp, 6'd0 };
assign lut_1_bit_7_fill = {lut_val_1_n_7_pp[13], lut_val_1_n_7_pp[13], lut_val_1_n_7_pp[13], lut_val_1_n_7_pp[13], lut_val_1_n_7_pp[13], lut_val_1_n_7_pp[13], lut_val_1_n_7_pp[13], lut_val_1_n_7_pp[13],  lut_val_1_n_7_pp, 7'd0 };
assign lut_1_bit_8_fill = {lut_val_1_n_8_pp[13], lut_val_1_n_8_pp[13], lut_val_1_n_8_pp[13], lut_val_1_n_8_pp[13], lut_val_1_n_8_pp[13], lut_val_1_n_8_pp[13], lut_val_1_n_8_pp[13],  lut_val_1_n_8_pp, 8'd0 };
assign lut_1_bit_9_fill = {lut_val_1_n_9_pp[13], lut_val_1_n_9_pp[13], lut_val_1_n_9_pp[13], lut_val_1_n_9_pp[13], lut_val_1_n_9_pp[13], lut_val_1_n_9_pp[13],  lut_val_1_n_9_pp, 9'd0 };
assign lut_1_bit_10_fill = {lut_val_1_n_10_pp[13], lut_val_1_n_10_pp[13], lut_val_1_n_10_pp[13], lut_val_1_n_10_pp[13], lut_val_1_n_10_pp[13],  lut_val_1_n_10_pp, 10'd0 };
assign lut_1_bit_11_fill = {lut_val_1_n_11_pp[13], lut_val_1_n_11_pp[13], lut_val_1_n_11_pp[13], lut_val_1_n_11_pp[13],  lut_val_1_n_11_pp, 11'd0 };
assign lut_1_bit_12_fill = {lut_val_1_n_12_pp[13], lut_val_1_n_12_pp[13], lut_val_1_n_12_pp[13],  lut_val_1_n_12_pp, 12'd0 };
assign lut_1_bit_13_fill = {lut_val_1_n_13_pp[13], lut_val_1_n_13_pp[13],  lut_val_1_n_13_pp, 13'd0 };
assign lut_1_bit_14_fill = {lut_val_1_n_14_pp[13],  lut_val_1_n_14_pp, 14'd0 };
assign lut_1_bit_15_fill = { lut_val_1_n_15_pp, 15'd0 };
wire [29:0] tree_1_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_0_fill), .bin(lut_1_bit_1_fill), .res(tree_1_pp_l_0_n_0_n) );
defparam Uadd_1_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_1_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_1_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_2_fill), .bin(lut_1_bit_3_fill), .res(tree_1_pp_l_0_n_1_n) );
defparam Uadd_1_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_1_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_1_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_4_fill), .bin(lut_1_bit_5_fill), .res(tree_1_pp_l_0_n_2_n) );
defparam Uadd_1_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_1_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_1_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_6_fill), .bin(lut_1_bit_7_fill), .res(tree_1_pp_l_0_n_3_n) );
defparam Uadd_1_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_1_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_1_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_8_fill), .bin(lut_1_bit_9_fill), .res(tree_1_pp_l_0_n_4_n) );
defparam Uadd_1_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_1_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_1_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_10_fill), .bin(lut_1_bit_11_fill), .res(tree_1_pp_l_0_n_5_n) );
defparam Uadd_1_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_1_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_1_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_12_fill), .bin(lut_1_bit_13_fill), .res(tree_1_pp_l_0_n_6_n) );
defparam Uadd_1_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_1_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_1_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_14_fill), .bin(lut_1_bit_15_fill), .res(tree_1_pp_l_0_n_7_n) );
defparam Uadd_1_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_1_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_1_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_1_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_0_n_0_n), .bin(tree_1_pp_l_0_n_1_n), .res(tree_1_pp_l_1_n_0_n) );
defparam Uadd_1_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_1_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_1_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_1_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_0_n_2_n), .bin(tree_1_pp_l_0_n_3_n), .res(tree_1_pp_l_1_n_1_n) );
defparam Uadd_1_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_1_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_1_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_1_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_0_n_4_n), .bin(tree_1_pp_l_0_n_5_n), .res(tree_1_pp_l_1_n_2_n) );
defparam Uadd_1_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_1_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_1_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_1_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_0_n_6_n), .bin(tree_1_pp_l_0_n_7_n), .res(tree_1_pp_l_1_n_3_n) );
defparam Uadd_1_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_1_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_1_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_1_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_1_n_0_n), .bin(tree_1_pp_l_1_n_1_n), .res(tree_1_pp_l_2_n_0_n) );
defparam Uadd_1_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_1_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_1_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_1_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_1_n_2_n), .bin(tree_1_pp_l_1_n_3_n), .res(tree_1_pp_l_2_n_1_n) );
defparam Uadd_1_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_1_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_1_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_1_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_2_n_0_n), .bin(tree_1_pp_l_2_n_1_n), .res(tree_1_pp_l_3_n_0_n) );
defparam Uadd_1_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_1_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_1_n;
assign lut_val_1_n=tree_1_pp_l_3_n_0_n;
wire [28:0] lut_2_bit_0_fill;
wire [28:0] lut_2_bit_1_fill;
wire [28:0] lut_2_bit_2_fill;
wire [28:0] lut_2_bit_3_fill;
wire [28:0] lut_2_bit_4_fill;
wire [28:0] lut_2_bit_5_fill;
wire [28:0] lut_2_bit_6_fill;
wire [28:0] lut_2_bit_7_fill;
wire [28:0] lut_2_bit_8_fill;
wire [28:0] lut_2_bit_9_fill;
wire [28:0] lut_2_bit_10_fill;
wire [28:0] lut_2_bit_11_fill;
wire [28:0] lut_2_bit_12_fill;
wire [28:0] lut_2_bit_13_fill;
wire [28:0] lut_2_bit_14_fill;
wire [28:0] lut_2_bit_15_fill;
assign lut_2_bit_0_fill = {lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13], lut_val_2_n_0_pp[13],  lut_val_2_n_0_pp };
assign lut_2_bit_1_fill = {lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13], lut_val_2_n_1_pp[13],  lut_val_2_n_1_pp, 1'd0 };
assign lut_2_bit_2_fill = {lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13], lut_val_2_n_2_pp[13],  lut_val_2_n_2_pp, 2'd0 };
assign lut_2_bit_3_fill = {lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13], lut_val_2_n_3_pp[13],  lut_val_2_n_3_pp, 3'd0 };
assign lut_2_bit_4_fill = {lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13], lut_val_2_n_4_pp[13],  lut_val_2_n_4_pp, 4'd0 };
assign lut_2_bit_5_fill = {lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13], lut_val_2_n_5_pp[13],  lut_val_2_n_5_pp, 5'd0 };
assign lut_2_bit_6_fill = {lut_val_2_n_6_pp[13], lut_val_2_n_6_pp[13], lut_val_2_n_6_pp[13], lut_val_2_n_6_pp[13], lut_val_2_n_6_pp[13], lut_val_2_n_6_pp[13], lut_val_2_n_6_pp[13], lut_val_2_n_6_pp[13], lut_val_2_n_6_pp[13],  lut_val_2_n_6_pp, 6'd0 };
assign lut_2_bit_7_fill = {lut_val_2_n_7_pp[13], lut_val_2_n_7_pp[13], lut_val_2_n_7_pp[13], lut_val_2_n_7_pp[13], lut_val_2_n_7_pp[13], lut_val_2_n_7_pp[13], lut_val_2_n_7_pp[13], lut_val_2_n_7_pp[13],  lut_val_2_n_7_pp, 7'd0 };
assign lut_2_bit_8_fill = {lut_val_2_n_8_pp[13], lut_val_2_n_8_pp[13], lut_val_2_n_8_pp[13], lut_val_2_n_8_pp[13], lut_val_2_n_8_pp[13], lut_val_2_n_8_pp[13], lut_val_2_n_8_pp[13],  lut_val_2_n_8_pp, 8'd0 };
assign lut_2_bit_9_fill = {lut_val_2_n_9_pp[13], lut_val_2_n_9_pp[13], lut_val_2_n_9_pp[13], lut_val_2_n_9_pp[13], lut_val_2_n_9_pp[13], lut_val_2_n_9_pp[13],  lut_val_2_n_9_pp, 9'd0 };
assign lut_2_bit_10_fill = {lut_val_2_n_10_pp[13], lut_val_2_n_10_pp[13], lut_val_2_n_10_pp[13], lut_val_2_n_10_pp[13], lut_val_2_n_10_pp[13],  lut_val_2_n_10_pp, 10'd0 };
assign lut_2_bit_11_fill = {lut_val_2_n_11_pp[13], lut_val_2_n_11_pp[13], lut_val_2_n_11_pp[13], lut_val_2_n_11_pp[13],  lut_val_2_n_11_pp, 11'd0 };
assign lut_2_bit_12_fill = {lut_val_2_n_12_pp[13], lut_val_2_n_12_pp[13], lut_val_2_n_12_pp[13],  lut_val_2_n_12_pp, 12'd0 };
assign lut_2_bit_13_fill = {lut_val_2_n_13_pp[13], lut_val_2_n_13_pp[13],  lut_val_2_n_13_pp, 13'd0 };
assign lut_2_bit_14_fill = {lut_val_2_n_14_pp[13],  lut_val_2_n_14_pp, 14'd0 };
assign lut_2_bit_15_fill = { lut_val_2_n_15_pp, 15'd0 };
wire [29:0] tree_2_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_0_fill), .bin(lut_2_bit_1_fill), .res(tree_2_pp_l_0_n_0_n) );
defparam Uadd_2_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_2_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_2_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_2_fill), .bin(lut_2_bit_3_fill), .res(tree_2_pp_l_0_n_1_n) );
defparam Uadd_2_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_2_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_2_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_4_fill), .bin(lut_2_bit_5_fill), .res(tree_2_pp_l_0_n_2_n) );
defparam Uadd_2_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_2_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_2_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_6_fill), .bin(lut_2_bit_7_fill), .res(tree_2_pp_l_0_n_3_n) );
defparam Uadd_2_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_2_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_2_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_8_fill), .bin(lut_2_bit_9_fill), .res(tree_2_pp_l_0_n_4_n) );
defparam Uadd_2_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_2_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_2_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_10_fill), .bin(lut_2_bit_11_fill), .res(tree_2_pp_l_0_n_5_n) );
defparam Uadd_2_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_2_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_2_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_12_fill), .bin(lut_2_bit_13_fill), .res(tree_2_pp_l_0_n_6_n) );
defparam Uadd_2_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_2_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_2_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_14_fill), .bin(lut_2_bit_15_fill), .res(tree_2_pp_l_0_n_7_n) );
defparam Uadd_2_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_2_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_2_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_2_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_0_n_0_n), .bin(tree_2_pp_l_0_n_1_n), .res(tree_2_pp_l_1_n_0_n) );
defparam Uadd_2_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_2_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_2_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_2_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_0_n_2_n), .bin(tree_2_pp_l_0_n_3_n), .res(tree_2_pp_l_1_n_1_n) );
defparam Uadd_2_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_2_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_2_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_2_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_0_n_4_n), .bin(tree_2_pp_l_0_n_5_n), .res(tree_2_pp_l_1_n_2_n) );
defparam Uadd_2_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_2_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_2_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_2_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_0_n_6_n), .bin(tree_2_pp_l_0_n_7_n), .res(tree_2_pp_l_1_n_3_n) );
defparam Uadd_2_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_2_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_2_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_2_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_1_n_0_n), .bin(tree_2_pp_l_1_n_1_n), .res(tree_2_pp_l_2_n_0_n) );
defparam Uadd_2_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_2_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_2_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_2_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_1_n_2_n), .bin(tree_2_pp_l_1_n_3_n), .res(tree_2_pp_l_2_n_1_n) );
defparam Uadd_2_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_2_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_2_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_2_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_2_n_0_n), .bin(tree_2_pp_l_2_n_1_n), .res(tree_2_pp_l_3_n_0_n) );
defparam Uadd_2_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_2_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_2_n;
assign lut_val_2_n=tree_2_pp_l_3_n_0_n;
wire [28:0] lut_3_bit_0_fill;
wire [28:0] lut_3_bit_1_fill;
wire [28:0] lut_3_bit_2_fill;
wire [28:0] lut_3_bit_3_fill;
wire [28:0] lut_3_bit_4_fill;
wire [28:0] lut_3_bit_5_fill;
wire [28:0] lut_3_bit_6_fill;
wire [28:0] lut_3_bit_7_fill;
wire [28:0] lut_3_bit_8_fill;
wire [28:0] lut_3_bit_9_fill;
wire [28:0] lut_3_bit_10_fill;
wire [28:0] lut_3_bit_11_fill;
wire [28:0] lut_3_bit_12_fill;
wire [28:0] lut_3_bit_13_fill;
wire [28:0] lut_3_bit_14_fill;
wire [28:0] lut_3_bit_15_fill;
assign lut_3_bit_0_fill = {lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13], lut_val_3_n_0_pp[13],  lut_val_3_n_0_pp };
assign lut_3_bit_1_fill = {lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13], lut_val_3_n_1_pp[13],  lut_val_3_n_1_pp, 1'd0 };
assign lut_3_bit_2_fill = {lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13], lut_val_3_n_2_pp[13],  lut_val_3_n_2_pp, 2'd0 };
assign lut_3_bit_3_fill = {lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13], lut_val_3_n_3_pp[13],  lut_val_3_n_3_pp, 3'd0 };
assign lut_3_bit_4_fill = {lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13], lut_val_3_n_4_pp[13],  lut_val_3_n_4_pp, 4'd0 };
assign lut_3_bit_5_fill = {lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13], lut_val_3_n_5_pp[13],  lut_val_3_n_5_pp, 5'd0 };
assign lut_3_bit_6_fill = {lut_val_3_n_6_pp[13], lut_val_3_n_6_pp[13], lut_val_3_n_6_pp[13], lut_val_3_n_6_pp[13], lut_val_3_n_6_pp[13], lut_val_3_n_6_pp[13], lut_val_3_n_6_pp[13], lut_val_3_n_6_pp[13], lut_val_3_n_6_pp[13],  lut_val_3_n_6_pp, 6'd0 };
assign lut_3_bit_7_fill = {lut_val_3_n_7_pp[13], lut_val_3_n_7_pp[13], lut_val_3_n_7_pp[13], lut_val_3_n_7_pp[13], lut_val_3_n_7_pp[13], lut_val_3_n_7_pp[13], lut_val_3_n_7_pp[13], lut_val_3_n_7_pp[13],  lut_val_3_n_7_pp, 7'd0 };
assign lut_3_bit_8_fill = {lut_val_3_n_8_pp[13], lut_val_3_n_8_pp[13], lut_val_3_n_8_pp[13], lut_val_3_n_8_pp[13], lut_val_3_n_8_pp[13], lut_val_3_n_8_pp[13], lut_val_3_n_8_pp[13],  lut_val_3_n_8_pp, 8'd0 };
assign lut_3_bit_9_fill = {lut_val_3_n_9_pp[13], lut_val_3_n_9_pp[13], lut_val_3_n_9_pp[13], lut_val_3_n_9_pp[13], lut_val_3_n_9_pp[13], lut_val_3_n_9_pp[13],  lut_val_3_n_9_pp, 9'd0 };
assign lut_3_bit_10_fill = {lut_val_3_n_10_pp[13], lut_val_3_n_10_pp[13], lut_val_3_n_10_pp[13], lut_val_3_n_10_pp[13], lut_val_3_n_10_pp[13],  lut_val_3_n_10_pp, 10'd0 };
assign lut_3_bit_11_fill = {lut_val_3_n_11_pp[13], lut_val_3_n_11_pp[13], lut_val_3_n_11_pp[13], lut_val_3_n_11_pp[13],  lut_val_3_n_11_pp, 11'd0 };
assign lut_3_bit_12_fill = {lut_val_3_n_12_pp[13], lut_val_3_n_12_pp[13], lut_val_3_n_12_pp[13],  lut_val_3_n_12_pp, 12'd0 };
assign lut_3_bit_13_fill = {lut_val_3_n_13_pp[13], lut_val_3_n_13_pp[13],  lut_val_3_n_13_pp, 13'd0 };
assign lut_3_bit_14_fill = {lut_val_3_n_14_pp[13],  lut_val_3_n_14_pp, 14'd0 };
assign lut_3_bit_15_fill = { lut_val_3_n_15_pp, 15'd0 };
wire [29:0] tree_3_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_0_fill), .bin(lut_3_bit_1_fill), .res(tree_3_pp_l_0_n_0_n) );
defparam Uadd_3_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_3_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_3_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_2_fill), .bin(lut_3_bit_3_fill), .res(tree_3_pp_l_0_n_1_n) );
defparam Uadd_3_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_3_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_3_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_4_fill), .bin(lut_3_bit_5_fill), .res(tree_3_pp_l_0_n_2_n) );
defparam Uadd_3_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_3_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_3_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_6_fill), .bin(lut_3_bit_7_fill), .res(tree_3_pp_l_0_n_3_n) );
defparam Uadd_3_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_3_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_3_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_8_fill), .bin(lut_3_bit_9_fill), .res(tree_3_pp_l_0_n_4_n) );
defparam Uadd_3_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_3_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_3_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_10_fill), .bin(lut_3_bit_11_fill), .res(tree_3_pp_l_0_n_5_n) );
defparam Uadd_3_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_3_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_3_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_12_fill), .bin(lut_3_bit_13_fill), .res(tree_3_pp_l_0_n_6_n) );
defparam Uadd_3_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_3_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_3_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_14_fill), .bin(lut_3_bit_15_fill), .res(tree_3_pp_l_0_n_7_n) );
defparam Uadd_3_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_3_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_3_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_3_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_0_n_0_n), .bin(tree_3_pp_l_0_n_1_n), .res(tree_3_pp_l_1_n_0_n) );
defparam Uadd_3_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_3_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_3_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_3_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_0_n_2_n), .bin(tree_3_pp_l_0_n_3_n), .res(tree_3_pp_l_1_n_1_n) );
defparam Uadd_3_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_3_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_3_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_3_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_0_n_4_n), .bin(tree_3_pp_l_0_n_5_n), .res(tree_3_pp_l_1_n_2_n) );
defparam Uadd_3_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_3_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_3_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_3_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_0_n_6_n), .bin(tree_3_pp_l_0_n_7_n), .res(tree_3_pp_l_1_n_3_n) );
defparam Uadd_3_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_3_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_3_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_3_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_1_n_0_n), .bin(tree_3_pp_l_1_n_1_n), .res(tree_3_pp_l_2_n_0_n) );
defparam Uadd_3_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_3_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_3_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_3_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_1_n_2_n), .bin(tree_3_pp_l_1_n_3_n), .res(tree_3_pp_l_2_n_1_n) );
defparam Uadd_3_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_3_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_3_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_3_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_2_n_0_n), .bin(tree_3_pp_l_2_n_1_n), .res(tree_3_pp_l_3_n_0_n) );
defparam Uadd_3_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_3_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_3_n;
assign lut_val_3_n=tree_3_pp_l_3_n_0_n;
wire [28:0] lut_4_bit_0_fill;
wire [28:0] lut_4_bit_1_fill;
wire [28:0] lut_4_bit_2_fill;
wire [28:0] lut_4_bit_3_fill;
wire [28:0] lut_4_bit_4_fill;
wire [28:0] lut_4_bit_5_fill;
wire [28:0] lut_4_bit_6_fill;
wire [28:0] lut_4_bit_7_fill;
wire [28:0] lut_4_bit_8_fill;
wire [28:0] lut_4_bit_9_fill;
wire [28:0] lut_4_bit_10_fill;
wire [28:0] lut_4_bit_11_fill;
wire [28:0] lut_4_bit_12_fill;
wire [28:0] lut_4_bit_13_fill;
wire [28:0] lut_4_bit_14_fill;
wire [28:0] lut_4_bit_15_fill;
assign lut_4_bit_0_fill = {lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13], lut_val_4_n_0_pp[13],  lut_val_4_n_0_pp };
assign lut_4_bit_1_fill = {lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13], lut_val_4_n_1_pp[13],  lut_val_4_n_1_pp, 1'd0 };
assign lut_4_bit_2_fill = {lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13], lut_val_4_n_2_pp[13],  lut_val_4_n_2_pp, 2'd0 };
assign lut_4_bit_3_fill = {lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13], lut_val_4_n_3_pp[13],  lut_val_4_n_3_pp, 3'd0 };
assign lut_4_bit_4_fill = {lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13], lut_val_4_n_4_pp[13],  lut_val_4_n_4_pp, 4'd0 };
assign lut_4_bit_5_fill = {lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13], lut_val_4_n_5_pp[13],  lut_val_4_n_5_pp, 5'd0 };
assign lut_4_bit_6_fill = {lut_val_4_n_6_pp[13], lut_val_4_n_6_pp[13], lut_val_4_n_6_pp[13], lut_val_4_n_6_pp[13], lut_val_4_n_6_pp[13], lut_val_4_n_6_pp[13], lut_val_4_n_6_pp[13], lut_val_4_n_6_pp[13], lut_val_4_n_6_pp[13],  lut_val_4_n_6_pp, 6'd0 };
assign lut_4_bit_7_fill = {lut_val_4_n_7_pp[13], lut_val_4_n_7_pp[13], lut_val_4_n_7_pp[13], lut_val_4_n_7_pp[13], lut_val_4_n_7_pp[13], lut_val_4_n_7_pp[13], lut_val_4_n_7_pp[13], lut_val_4_n_7_pp[13],  lut_val_4_n_7_pp, 7'd0 };
assign lut_4_bit_8_fill = {lut_val_4_n_8_pp[13], lut_val_4_n_8_pp[13], lut_val_4_n_8_pp[13], lut_val_4_n_8_pp[13], lut_val_4_n_8_pp[13], lut_val_4_n_8_pp[13], lut_val_4_n_8_pp[13],  lut_val_4_n_8_pp, 8'd0 };
assign lut_4_bit_9_fill = {lut_val_4_n_9_pp[13], lut_val_4_n_9_pp[13], lut_val_4_n_9_pp[13], lut_val_4_n_9_pp[13], lut_val_4_n_9_pp[13], lut_val_4_n_9_pp[13],  lut_val_4_n_9_pp, 9'd0 };
assign lut_4_bit_10_fill = {lut_val_4_n_10_pp[13], lut_val_4_n_10_pp[13], lut_val_4_n_10_pp[13], lut_val_4_n_10_pp[13], lut_val_4_n_10_pp[13],  lut_val_4_n_10_pp, 10'd0 };
assign lut_4_bit_11_fill = {lut_val_4_n_11_pp[13], lut_val_4_n_11_pp[13], lut_val_4_n_11_pp[13], lut_val_4_n_11_pp[13],  lut_val_4_n_11_pp, 11'd0 };
assign lut_4_bit_12_fill = {lut_val_4_n_12_pp[13], lut_val_4_n_12_pp[13], lut_val_4_n_12_pp[13],  lut_val_4_n_12_pp, 12'd0 };
assign lut_4_bit_13_fill = {lut_val_4_n_13_pp[13], lut_val_4_n_13_pp[13],  lut_val_4_n_13_pp, 13'd0 };
assign lut_4_bit_14_fill = {lut_val_4_n_14_pp[13],  lut_val_4_n_14_pp, 14'd0 };
assign lut_4_bit_15_fill = { lut_val_4_n_15_pp, 15'd0 };
wire [29:0] tree_4_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_4_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_4_bit_0_fill), .bin(lut_4_bit_1_fill), .res(tree_4_pp_l_0_n_0_n) );
defparam Uadd_4_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_4_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_4_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_4_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_4_bit_2_fill), .bin(lut_4_bit_3_fill), .res(tree_4_pp_l_0_n_1_n) );
defparam Uadd_4_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_4_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_4_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_4_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_4_bit_4_fill), .bin(lut_4_bit_5_fill), .res(tree_4_pp_l_0_n_2_n) );
defparam Uadd_4_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_4_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_4_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_4_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_4_bit_6_fill), .bin(lut_4_bit_7_fill), .res(tree_4_pp_l_0_n_3_n) );
defparam Uadd_4_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_4_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_4_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_4_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_4_bit_8_fill), .bin(lut_4_bit_9_fill), .res(tree_4_pp_l_0_n_4_n) );
defparam Uadd_4_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_4_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_4_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_4_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_4_bit_10_fill), .bin(lut_4_bit_11_fill), .res(tree_4_pp_l_0_n_5_n) );
defparam Uadd_4_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_4_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_4_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_4_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_4_bit_12_fill), .bin(lut_4_bit_13_fill), .res(tree_4_pp_l_0_n_6_n) );
defparam Uadd_4_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_4_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_4_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_4_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_4_bit_14_fill), .bin(lut_4_bit_15_fill), .res(tree_4_pp_l_0_n_7_n) );
defparam Uadd_4_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_4_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_4_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_4_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_4_pp_l_0_n_0_n), .bin(tree_4_pp_l_0_n_1_n), .res(tree_4_pp_l_1_n_0_n) );
defparam Uadd_4_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_4_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_4_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_4_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_4_pp_l_0_n_2_n), .bin(tree_4_pp_l_0_n_3_n), .res(tree_4_pp_l_1_n_1_n) );
defparam Uadd_4_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_4_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_4_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_4_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_4_pp_l_0_n_4_n), .bin(tree_4_pp_l_0_n_5_n), .res(tree_4_pp_l_1_n_2_n) );
defparam Uadd_4_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_4_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_4_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_4_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_4_pp_l_0_n_6_n), .bin(tree_4_pp_l_0_n_7_n), .res(tree_4_pp_l_1_n_3_n) );
defparam Uadd_4_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_4_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_4_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_4_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_4_pp_l_1_n_0_n), .bin(tree_4_pp_l_1_n_1_n), .res(tree_4_pp_l_2_n_0_n) );
defparam Uadd_4_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_4_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_4_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_4_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_4_pp_l_1_n_2_n), .bin(tree_4_pp_l_1_n_3_n), .res(tree_4_pp_l_2_n_1_n) );
defparam Uadd_4_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_4_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_4_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_4_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_4_pp_l_2_n_0_n), .bin(tree_4_pp_l_2_n_1_n), .res(tree_4_pp_l_3_n_0_n) );
defparam Uadd_4_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_4_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_4_n;
assign lut_val_4_n=tree_4_pp_l_3_n_0_n;
wire [28:0] lut_5_bit_0_fill;
wire [28:0] lut_5_bit_1_fill;
wire [28:0] lut_5_bit_2_fill;
wire [28:0] lut_5_bit_3_fill;
wire [28:0] lut_5_bit_4_fill;
wire [28:0] lut_5_bit_5_fill;
wire [28:0] lut_5_bit_6_fill;
wire [28:0] lut_5_bit_7_fill;
wire [28:0] lut_5_bit_8_fill;
wire [28:0] lut_5_bit_9_fill;
wire [28:0] lut_5_bit_10_fill;
wire [28:0] lut_5_bit_11_fill;
wire [28:0] lut_5_bit_12_fill;
wire [28:0] lut_5_bit_13_fill;
wire [28:0] lut_5_bit_14_fill;
wire [28:0] lut_5_bit_15_fill;
assign lut_5_bit_0_fill = {lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13], lut_val_5_n_0_pp[13],  lut_val_5_n_0_pp };
assign lut_5_bit_1_fill = {lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13], lut_val_5_n_1_pp[13],  lut_val_5_n_1_pp, 1'd0 };
assign lut_5_bit_2_fill = {lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13], lut_val_5_n_2_pp[13],  lut_val_5_n_2_pp, 2'd0 };
assign lut_5_bit_3_fill = {lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13], lut_val_5_n_3_pp[13],  lut_val_5_n_3_pp, 3'd0 };
assign lut_5_bit_4_fill = {lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13], lut_val_5_n_4_pp[13],  lut_val_5_n_4_pp, 4'd0 };
assign lut_5_bit_5_fill = {lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13], lut_val_5_n_5_pp[13],  lut_val_5_n_5_pp, 5'd0 };
assign lut_5_bit_6_fill = {lut_val_5_n_6_pp[13], lut_val_5_n_6_pp[13], lut_val_5_n_6_pp[13], lut_val_5_n_6_pp[13], lut_val_5_n_6_pp[13], lut_val_5_n_6_pp[13], lut_val_5_n_6_pp[13], lut_val_5_n_6_pp[13], lut_val_5_n_6_pp[13],  lut_val_5_n_6_pp, 6'd0 };
assign lut_5_bit_7_fill = {lut_val_5_n_7_pp[13], lut_val_5_n_7_pp[13], lut_val_5_n_7_pp[13], lut_val_5_n_7_pp[13], lut_val_5_n_7_pp[13], lut_val_5_n_7_pp[13], lut_val_5_n_7_pp[13], lut_val_5_n_7_pp[13],  lut_val_5_n_7_pp, 7'd0 };
assign lut_5_bit_8_fill = {lut_val_5_n_8_pp[13], lut_val_5_n_8_pp[13], lut_val_5_n_8_pp[13], lut_val_5_n_8_pp[13], lut_val_5_n_8_pp[13], lut_val_5_n_8_pp[13], lut_val_5_n_8_pp[13],  lut_val_5_n_8_pp, 8'd0 };
assign lut_5_bit_9_fill = {lut_val_5_n_9_pp[13], lut_val_5_n_9_pp[13], lut_val_5_n_9_pp[13], lut_val_5_n_9_pp[13], lut_val_5_n_9_pp[13], lut_val_5_n_9_pp[13],  lut_val_5_n_9_pp, 9'd0 };
assign lut_5_bit_10_fill = {lut_val_5_n_10_pp[13], lut_val_5_n_10_pp[13], lut_val_5_n_10_pp[13], lut_val_5_n_10_pp[13], lut_val_5_n_10_pp[13],  lut_val_5_n_10_pp, 10'd0 };
assign lut_5_bit_11_fill = {lut_val_5_n_11_pp[13], lut_val_5_n_11_pp[13], lut_val_5_n_11_pp[13], lut_val_5_n_11_pp[13],  lut_val_5_n_11_pp, 11'd0 };
assign lut_5_bit_12_fill = {lut_val_5_n_12_pp[13], lut_val_5_n_12_pp[13], lut_val_5_n_12_pp[13],  lut_val_5_n_12_pp, 12'd0 };
assign lut_5_bit_13_fill = {lut_val_5_n_13_pp[13], lut_val_5_n_13_pp[13],  lut_val_5_n_13_pp, 13'd0 };
assign lut_5_bit_14_fill = {lut_val_5_n_14_pp[13],  lut_val_5_n_14_pp, 14'd0 };
assign lut_5_bit_15_fill = { lut_val_5_n_15_pp, 15'd0 };
wire [29:0] tree_5_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_5_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_5_bit_0_fill), .bin(lut_5_bit_1_fill), .res(tree_5_pp_l_0_n_0_n) );
defparam Uadd_5_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_5_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_5_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_5_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_5_bit_2_fill), .bin(lut_5_bit_3_fill), .res(tree_5_pp_l_0_n_1_n) );
defparam Uadd_5_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_5_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_5_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_5_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_5_bit_4_fill), .bin(lut_5_bit_5_fill), .res(tree_5_pp_l_0_n_2_n) );
defparam Uadd_5_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_5_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_5_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_5_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_5_bit_6_fill), .bin(lut_5_bit_7_fill), .res(tree_5_pp_l_0_n_3_n) );
defparam Uadd_5_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_5_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_5_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_5_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_5_bit_8_fill), .bin(lut_5_bit_9_fill), .res(tree_5_pp_l_0_n_4_n) );
defparam Uadd_5_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_5_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_5_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_5_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_5_bit_10_fill), .bin(lut_5_bit_11_fill), .res(tree_5_pp_l_0_n_5_n) );
defparam Uadd_5_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_5_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_5_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_5_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_5_bit_12_fill), .bin(lut_5_bit_13_fill), .res(tree_5_pp_l_0_n_6_n) );
defparam Uadd_5_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_5_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_5_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_5_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_5_bit_14_fill), .bin(lut_5_bit_15_fill), .res(tree_5_pp_l_0_n_7_n) );
defparam Uadd_5_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_5_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_5_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_5_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_5_pp_l_0_n_0_n), .bin(tree_5_pp_l_0_n_1_n), .res(tree_5_pp_l_1_n_0_n) );
defparam Uadd_5_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_5_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_5_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_5_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_5_pp_l_0_n_2_n), .bin(tree_5_pp_l_0_n_3_n), .res(tree_5_pp_l_1_n_1_n) );
defparam Uadd_5_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_5_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_5_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_5_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_5_pp_l_0_n_4_n), .bin(tree_5_pp_l_0_n_5_n), .res(tree_5_pp_l_1_n_2_n) );
defparam Uadd_5_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_5_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_5_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_5_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_5_pp_l_0_n_6_n), .bin(tree_5_pp_l_0_n_7_n), .res(tree_5_pp_l_1_n_3_n) );
defparam Uadd_5_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_5_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_5_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_5_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_5_pp_l_1_n_0_n), .bin(tree_5_pp_l_1_n_1_n), .res(tree_5_pp_l_2_n_0_n) );
defparam Uadd_5_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_5_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_5_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_5_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_5_pp_l_1_n_2_n), .bin(tree_5_pp_l_1_n_3_n), .res(tree_5_pp_l_2_n_1_n) );
defparam Uadd_5_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_5_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_5_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_5_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_5_pp_l_2_n_0_n), .bin(tree_5_pp_l_2_n_1_n), .res(tree_5_pp_l_3_n_0_n) );
defparam Uadd_5_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_5_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_5_n;
assign lut_val_5_n=tree_5_pp_l_3_n_0_n;
wire [28:0] lut_6_bit_0_fill;
wire [28:0] lut_6_bit_1_fill;
wire [28:0] lut_6_bit_2_fill;
wire [28:0] lut_6_bit_3_fill;
wire [28:0] lut_6_bit_4_fill;
wire [28:0] lut_6_bit_5_fill;
wire [28:0] lut_6_bit_6_fill;
wire [28:0] lut_6_bit_7_fill;
wire [28:0] lut_6_bit_8_fill;
wire [28:0] lut_6_bit_9_fill;
wire [28:0] lut_6_bit_10_fill;
wire [28:0] lut_6_bit_11_fill;
wire [28:0] lut_6_bit_12_fill;
wire [28:0] lut_6_bit_13_fill;
wire [28:0] lut_6_bit_14_fill;
wire [28:0] lut_6_bit_15_fill;
assign lut_6_bit_0_fill = {lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13], lut_val_6_n_0_pp[13],  lut_val_6_n_0_pp };
assign lut_6_bit_1_fill = {lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13], lut_val_6_n_1_pp[13],  lut_val_6_n_1_pp, 1'd0 };
assign lut_6_bit_2_fill = {lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13], lut_val_6_n_2_pp[13],  lut_val_6_n_2_pp, 2'd0 };
assign lut_6_bit_3_fill = {lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13], lut_val_6_n_3_pp[13],  lut_val_6_n_3_pp, 3'd0 };
assign lut_6_bit_4_fill = {lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13], lut_val_6_n_4_pp[13],  lut_val_6_n_4_pp, 4'd0 };
assign lut_6_bit_5_fill = {lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13], lut_val_6_n_5_pp[13],  lut_val_6_n_5_pp, 5'd0 };
assign lut_6_bit_6_fill = {lut_val_6_n_6_pp[13], lut_val_6_n_6_pp[13], lut_val_6_n_6_pp[13], lut_val_6_n_6_pp[13], lut_val_6_n_6_pp[13], lut_val_6_n_6_pp[13], lut_val_6_n_6_pp[13], lut_val_6_n_6_pp[13], lut_val_6_n_6_pp[13],  lut_val_6_n_6_pp, 6'd0 };
assign lut_6_bit_7_fill = {lut_val_6_n_7_pp[13], lut_val_6_n_7_pp[13], lut_val_6_n_7_pp[13], lut_val_6_n_7_pp[13], lut_val_6_n_7_pp[13], lut_val_6_n_7_pp[13], lut_val_6_n_7_pp[13], lut_val_6_n_7_pp[13],  lut_val_6_n_7_pp, 7'd0 };
assign lut_6_bit_8_fill = {lut_val_6_n_8_pp[13], lut_val_6_n_8_pp[13], lut_val_6_n_8_pp[13], lut_val_6_n_8_pp[13], lut_val_6_n_8_pp[13], lut_val_6_n_8_pp[13], lut_val_6_n_8_pp[13],  lut_val_6_n_8_pp, 8'd0 };
assign lut_6_bit_9_fill = {lut_val_6_n_9_pp[13], lut_val_6_n_9_pp[13], lut_val_6_n_9_pp[13], lut_val_6_n_9_pp[13], lut_val_6_n_9_pp[13], lut_val_6_n_9_pp[13],  lut_val_6_n_9_pp, 9'd0 };
assign lut_6_bit_10_fill = {lut_val_6_n_10_pp[13], lut_val_6_n_10_pp[13], lut_val_6_n_10_pp[13], lut_val_6_n_10_pp[13], lut_val_6_n_10_pp[13],  lut_val_6_n_10_pp, 10'd0 };
assign lut_6_bit_11_fill = {lut_val_6_n_11_pp[13], lut_val_6_n_11_pp[13], lut_val_6_n_11_pp[13], lut_val_6_n_11_pp[13],  lut_val_6_n_11_pp, 11'd0 };
assign lut_6_bit_12_fill = {lut_val_6_n_12_pp[13], lut_val_6_n_12_pp[13], lut_val_6_n_12_pp[13],  lut_val_6_n_12_pp, 12'd0 };
assign lut_6_bit_13_fill = {lut_val_6_n_13_pp[13], lut_val_6_n_13_pp[13],  lut_val_6_n_13_pp, 13'd0 };
assign lut_6_bit_14_fill = {lut_val_6_n_14_pp[13],  lut_val_6_n_14_pp, 14'd0 };
assign lut_6_bit_15_fill = { lut_val_6_n_15_pp, 15'd0 };
wire [29:0] tree_6_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_6_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_6_bit_0_fill), .bin(lut_6_bit_1_fill), .res(tree_6_pp_l_0_n_0_n) );
defparam Uadd_6_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_6_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_6_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_6_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_6_bit_2_fill), .bin(lut_6_bit_3_fill), .res(tree_6_pp_l_0_n_1_n) );
defparam Uadd_6_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_6_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_6_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_6_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_6_bit_4_fill), .bin(lut_6_bit_5_fill), .res(tree_6_pp_l_0_n_2_n) );
defparam Uadd_6_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_6_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_6_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_6_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_6_bit_6_fill), .bin(lut_6_bit_7_fill), .res(tree_6_pp_l_0_n_3_n) );
defparam Uadd_6_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_6_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_6_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_6_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_6_bit_8_fill), .bin(lut_6_bit_9_fill), .res(tree_6_pp_l_0_n_4_n) );
defparam Uadd_6_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_6_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_6_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_6_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_6_bit_10_fill), .bin(lut_6_bit_11_fill), .res(tree_6_pp_l_0_n_5_n) );
defparam Uadd_6_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_6_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_6_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_6_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_6_bit_12_fill), .bin(lut_6_bit_13_fill), .res(tree_6_pp_l_0_n_6_n) );
defparam Uadd_6_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_6_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_6_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_6_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_6_bit_14_fill), .bin(lut_6_bit_15_fill), .res(tree_6_pp_l_0_n_7_n) );
defparam Uadd_6_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_6_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_6_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_6_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_6_pp_l_0_n_0_n), .bin(tree_6_pp_l_0_n_1_n), .res(tree_6_pp_l_1_n_0_n) );
defparam Uadd_6_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_6_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_6_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_6_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_6_pp_l_0_n_2_n), .bin(tree_6_pp_l_0_n_3_n), .res(tree_6_pp_l_1_n_1_n) );
defparam Uadd_6_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_6_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_6_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_6_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_6_pp_l_0_n_4_n), .bin(tree_6_pp_l_0_n_5_n), .res(tree_6_pp_l_1_n_2_n) );
defparam Uadd_6_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_6_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_6_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_6_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_6_pp_l_0_n_6_n), .bin(tree_6_pp_l_0_n_7_n), .res(tree_6_pp_l_1_n_3_n) );
defparam Uadd_6_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_6_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_6_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_6_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_6_pp_l_1_n_0_n), .bin(tree_6_pp_l_1_n_1_n), .res(tree_6_pp_l_2_n_0_n) );
defparam Uadd_6_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_6_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_6_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_6_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_6_pp_l_1_n_2_n), .bin(tree_6_pp_l_1_n_3_n), .res(tree_6_pp_l_2_n_1_n) );
defparam Uadd_6_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_6_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_6_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_6_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_6_pp_l_2_n_0_n), .bin(tree_6_pp_l_2_n_1_n), .res(tree_6_pp_l_3_n_0_n) );
defparam Uadd_6_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_6_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_6_n;
assign lut_val_6_n=tree_6_pp_l_3_n_0_n;
wire [28:0] lut_7_bit_0_fill;
wire [28:0] lut_7_bit_1_fill;
wire [28:0] lut_7_bit_2_fill;
wire [28:0] lut_7_bit_3_fill;
wire [28:0] lut_7_bit_4_fill;
wire [28:0] lut_7_bit_5_fill;
wire [28:0] lut_7_bit_6_fill;
wire [28:0] lut_7_bit_7_fill;
wire [28:0] lut_7_bit_8_fill;
wire [28:0] lut_7_bit_9_fill;
wire [28:0] lut_7_bit_10_fill;
wire [28:0] lut_7_bit_11_fill;
wire [28:0] lut_7_bit_12_fill;
wire [28:0] lut_7_bit_13_fill;
wire [28:0] lut_7_bit_14_fill;
wire [28:0] lut_7_bit_15_fill;
assign lut_7_bit_0_fill = {lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13], lut_val_7_n_0_pp[13],  lut_val_7_n_0_pp };
assign lut_7_bit_1_fill = {lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13], lut_val_7_n_1_pp[13],  lut_val_7_n_1_pp, 1'd0 };
assign lut_7_bit_2_fill = {lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13], lut_val_7_n_2_pp[13],  lut_val_7_n_2_pp, 2'd0 };
assign lut_7_bit_3_fill = {lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13], lut_val_7_n_3_pp[13],  lut_val_7_n_3_pp, 3'd0 };
assign lut_7_bit_4_fill = {lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13], lut_val_7_n_4_pp[13],  lut_val_7_n_4_pp, 4'd0 };
assign lut_7_bit_5_fill = {lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13], lut_val_7_n_5_pp[13],  lut_val_7_n_5_pp, 5'd0 };
assign lut_7_bit_6_fill = {lut_val_7_n_6_pp[13], lut_val_7_n_6_pp[13], lut_val_7_n_6_pp[13], lut_val_7_n_6_pp[13], lut_val_7_n_6_pp[13], lut_val_7_n_6_pp[13], lut_val_7_n_6_pp[13], lut_val_7_n_6_pp[13], lut_val_7_n_6_pp[13],  lut_val_7_n_6_pp, 6'd0 };
assign lut_7_bit_7_fill = {lut_val_7_n_7_pp[13], lut_val_7_n_7_pp[13], lut_val_7_n_7_pp[13], lut_val_7_n_7_pp[13], lut_val_7_n_7_pp[13], lut_val_7_n_7_pp[13], lut_val_7_n_7_pp[13], lut_val_7_n_7_pp[13],  lut_val_7_n_7_pp, 7'd0 };
assign lut_7_bit_8_fill = {lut_val_7_n_8_pp[13], lut_val_7_n_8_pp[13], lut_val_7_n_8_pp[13], lut_val_7_n_8_pp[13], lut_val_7_n_8_pp[13], lut_val_7_n_8_pp[13], lut_val_7_n_8_pp[13],  lut_val_7_n_8_pp, 8'd0 };
assign lut_7_bit_9_fill = {lut_val_7_n_9_pp[13], lut_val_7_n_9_pp[13], lut_val_7_n_9_pp[13], lut_val_7_n_9_pp[13], lut_val_7_n_9_pp[13], lut_val_7_n_9_pp[13],  lut_val_7_n_9_pp, 9'd0 };
assign lut_7_bit_10_fill = {lut_val_7_n_10_pp[13], lut_val_7_n_10_pp[13], lut_val_7_n_10_pp[13], lut_val_7_n_10_pp[13], lut_val_7_n_10_pp[13],  lut_val_7_n_10_pp, 10'd0 };
assign lut_7_bit_11_fill = {lut_val_7_n_11_pp[13], lut_val_7_n_11_pp[13], lut_val_7_n_11_pp[13], lut_val_7_n_11_pp[13],  lut_val_7_n_11_pp, 11'd0 };
assign lut_7_bit_12_fill = {lut_val_7_n_12_pp[13], lut_val_7_n_12_pp[13], lut_val_7_n_12_pp[13],  lut_val_7_n_12_pp, 12'd0 };
assign lut_7_bit_13_fill = {lut_val_7_n_13_pp[13], lut_val_7_n_13_pp[13],  lut_val_7_n_13_pp, 13'd0 };
assign lut_7_bit_14_fill = {lut_val_7_n_14_pp[13],  lut_val_7_n_14_pp, 14'd0 };
assign lut_7_bit_15_fill = { lut_val_7_n_15_pp, 15'd0 };
wire [29:0] tree_7_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_7_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_7_bit_0_fill), .bin(lut_7_bit_1_fill), .res(tree_7_pp_l_0_n_0_n) );
defparam Uadd_7_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_7_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_7_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_7_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_7_bit_2_fill), .bin(lut_7_bit_3_fill), .res(tree_7_pp_l_0_n_1_n) );
defparam Uadd_7_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_7_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_7_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_7_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_7_bit_4_fill), .bin(lut_7_bit_5_fill), .res(tree_7_pp_l_0_n_2_n) );
defparam Uadd_7_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_7_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_7_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_7_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_7_bit_6_fill), .bin(lut_7_bit_7_fill), .res(tree_7_pp_l_0_n_3_n) );
defparam Uadd_7_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_7_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_7_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_7_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_7_bit_8_fill), .bin(lut_7_bit_9_fill), .res(tree_7_pp_l_0_n_4_n) );
defparam Uadd_7_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_7_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_7_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_7_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_7_bit_10_fill), .bin(lut_7_bit_11_fill), .res(tree_7_pp_l_0_n_5_n) );
defparam Uadd_7_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_7_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_7_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_7_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_7_bit_12_fill), .bin(lut_7_bit_13_fill), .res(tree_7_pp_l_0_n_6_n) );
defparam Uadd_7_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_7_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_7_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_7_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_7_bit_14_fill), .bin(lut_7_bit_15_fill), .res(tree_7_pp_l_0_n_7_n) );
defparam Uadd_7_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_7_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_7_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_7_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_7_pp_l_0_n_0_n), .bin(tree_7_pp_l_0_n_1_n), .res(tree_7_pp_l_1_n_0_n) );
defparam Uadd_7_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_7_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_7_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_7_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_7_pp_l_0_n_2_n), .bin(tree_7_pp_l_0_n_3_n), .res(tree_7_pp_l_1_n_1_n) );
defparam Uadd_7_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_7_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_7_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_7_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_7_pp_l_0_n_4_n), .bin(tree_7_pp_l_0_n_5_n), .res(tree_7_pp_l_1_n_2_n) );
defparam Uadd_7_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_7_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_7_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_7_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_7_pp_l_0_n_6_n), .bin(tree_7_pp_l_0_n_7_n), .res(tree_7_pp_l_1_n_3_n) );
defparam Uadd_7_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_7_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_7_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_7_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_7_pp_l_1_n_0_n), .bin(tree_7_pp_l_1_n_1_n), .res(tree_7_pp_l_2_n_0_n) );
defparam Uadd_7_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_7_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_7_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_7_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_7_pp_l_1_n_2_n), .bin(tree_7_pp_l_1_n_3_n), .res(tree_7_pp_l_2_n_1_n) );
defparam Uadd_7_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_7_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_7_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_7_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_7_pp_l_2_n_0_n), .bin(tree_7_pp_l_2_n_1_n), .res(tree_7_pp_l_3_n_0_n) );
defparam Uadd_7_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_7_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_7_n;
assign lut_val_7_n=tree_7_pp_l_3_n_0_n;
wire [28:0] lut_8_bit_0_fill;
wire [28:0] lut_8_bit_1_fill;
wire [28:0] lut_8_bit_2_fill;
wire [28:0] lut_8_bit_3_fill;
wire [28:0] lut_8_bit_4_fill;
wire [28:0] lut_8_bit_5_fill;
wire [28:0] lut_8_bit_6_fill;
wire [28:0] lut_8_bit_7_fill;
wire [28:0] lut_8_bit_8_fill;
wire [28:0] lut_8_bit_9_fill;
wire [28:0] lut_8_bit_10_fill;
wire [28:0] lut_8_bit_11_fill;
wire [28:0] lut_8_bit_12_fill;
wire [28:0] lut_8_bit_13_fill;
wire [28:0] lut_8_bit_14_fill;
wire [28:0] lut_8_bit_15_fill;
assign lut_8_bit_0_fill = {lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13], lut_val_8_n_0_pp[13],  lut_val_8_n_0_pp };
assign lut_8_bit_1_fill = {lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13], lut_val_8_n_1_pp[13],  lut_val_8_n_1_pp, 1'd0 };
assign lut_8_bit_2_fill = {lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13], lut_val_8_n_2_pp[13],  lut_val_8_n_2_pp, 2'd0 };
assign lut_8_bit_3_fill = {lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13], lut_val_8_n_3_pp[13],  lut_val_8_n_3_pp, 3'd0 };
assign lut_8_bit_4_fill = {lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13], lut_val_8_n_4_pp[13],  lut_val_8_n_4_pp, 4'd0 };
assign lut_8_bit_5_fill = {lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13], lut_val_8_n_5_pp[13],  lut_val_8_n_5_pp, 5'd0 };
assign lut_8_bit_6_fill = {lut_val_8_n_6_pp[13], lut_val_8_n_6_pp[13], lut_val_8_n_6_pp[13], lut_val_8_n_6_pp[13], lut_val_8_n_6_pp[13], lut_val_8_n_6_pp[13], lut_val_8_n_6_pp[13], lut_val_8_n_6_pp[13], lut_val_8_n_6_pp[13],  lut_val_8_n_6_pp, 6'd0 };
assign lut_8_bit_7_fill = {lut_val_8_n_7_pp[13], lut_val_8_n_7_pp[13], lut_val_8_n_7_pp[13], lut_val_8_n_7_pp[13], lut_val_8_n_7_pp[13], lut_val_8_n_7_pp[13], lut_val_8_n_7_pp[13], lut_val_8_n_7_pp[13],  lut_val_8_n_7_pp, 7'd0 };
assign lut_8_bit_8_fill = {lut_val_8_n_8_pp[13], lut_val_8_n_8_pp[13], lut_val_8_n_8_pp[13], lut_val_8_n_8_pp[13], lut_val_8_n_8_pp[13], lut_val_8_n_8_pp[13], lut_val_8_n_8_pp[13],  lut_val_8_n_8_pp, 8'd0 };
assign lut_8_bit_9_fill = {lut_val_8_n_9_pp[13], lut_val_8_n_9_pp[13], lut_val_8_n_9_pp[13], lut_val_8_n_9_pp[13], lut_val_8_n_9_pp[13], lut_val_8_n_9_pp[13],  lut_val_8_n_9_pp, 9'd0 };
assign lut_8_bit_10_fill = {lut_val_8_n_10_pp[13], lut_val_8_n_10_pp[13], lut_val_8_n_10_pp[13], lut_val_8_n_10_pp[13], lut_val_8_n_10_pp[13],  lut_val_8_n_10_pp, 10'd0 };
assign lut_8_bit_11_fill = {lut_val_8_n_11_pp[13], lut_val_8_n_11_pp[13], lut_val_8_n_11_pp[13], lut_val_8_n_11_pp[13],  lut_val_8_n_11_pp, 11'd0 };
assign lut_8_bit_12_fill = {lut_val_8_n_12_pp[13], lut_val_8_n_12_pp[13], lut_val_8_n_12_pp[13],  lut_val_8_n_12_pp, 12'd0 };
assign lut_8_bit_13_fill = {lut_val_8_n_13_pp[13], lut_val_8_n_13_pp[13],  lut_val_8_n_13_pp, 13'd0 };
assign lut_8_bit_14_fill = {lut_val_8_n_14_pp[13],  lut_val_8_n_14_pp, 14'd0 };
assign lut_8_bit_15_fill = { lut_val_8_n_15_pp, 15'd0 };
wire [29:0] tree_8_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_8_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_8_bit_0_fill), .bin(lut_8_bit_1_fill), .res(tree_8_pp_l_0_n_0_n) );
defparam Uadd_8_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_8_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_8_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_8_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_8_bit_2_fill), .bin(lut_8_bit_3_fill), .res(tree_8_pp_l_0_n_1_n) );
defparam Uadd_8_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_8_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_8_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_8_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_8_bit_4_fill), .bin(lut_8_bit_5_fill), .res(tree_8_pp_l_0_n_2_n) );
defparam Uadd_8_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_8_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_8_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_8_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_8_bit_6_fill), .bin(lut_8_bit_7_fill), .res(tree_8_pp_l_0_n_3_n) );
defparam Uadd_8_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_8_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_8_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_8_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_8_bit_8_fill), .bin(lut_8_bit_9_fill), .res(tree_8_pp_l_0_n_4_n) );
defparam Uadd_8_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_8_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_8_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_8_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_8_bit_10_fill), .bin(lut_8_bit_11_fill), .res(tree_8_pp_l_0_n_5_n) );
defparam Uadd_8_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_8_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_8_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_8_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_8_bit_12_fill), .bin(lut_8_bit_13_fill), .res(tree_8_pp_l_0_n_6_n) );
defparam Uadd_8_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_8_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_8_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_8_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_8_bit_14_fill), .bin(lut_8_bit_15_fill), .res(tree_8_pp_l_0_n_7_n) );
defparam Uadd_8_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_8_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_8_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_8_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_8_pp_l_0_n_0_n), .bin(tree_8_pp_l_0_n_1_n), .res(tree_8_pp_l_1_n_0_n) );
defparam Uadd_8_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_8_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_8_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_8_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_8_pp_l_0_n_2_n), .bin(tree_8_pp_l_0_n_3_n), .res(tree_8_pp_l_1_n_1_n) );
defparam Uadd_8_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_8_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_8_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_8_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_8_pp_l_0_n_4_n), .bin(tree_8_pp_l_0_n_5_n), .res(tree_8_pp_l_1_n_2_n) );
defparam Uadd_8_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_8_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_8_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_8_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_8_pp_l_0_n_6_n), .bin(tree_8_pp_l_0_n_7_n), .res(tree_8_pp_l_1_n_3_n) );
defparam Uadd_8_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_8_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_8_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_8_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_8_pp_l_1_n_0_n), .bin(tree_8_pp_l_1_n_1_n), .res(tree_8_pp_l_2_n_0_n) );
defparam Uadd_8_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_8_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_8_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_8_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_8_pp_l_1_n_2_n), .bin(tree_8_pp_l_1_n_3_n), .res(tree_8_pp_l_2_n_1_n) );
defparam Uadd_8_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_8_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_8_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_8_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_8_pp_l_2_n_0_n), .bin(tree_8_pp_l_2_n_1_n), .res(tree_8_pp_l_3_n_0_n) );
defparam Uadd_8_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_8_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_8_n;
assign lut_val_8_n=tree_8_pp_l_3_n_0_n;
wire [28:0] lut_9_bit_0_fill;
wire [28:0] lut_9_bit_1_fill;
wire [28:0] lut_9_bit_2_fill;
wire [28:0] lut_9_bit_3_fill;
wire [28:0] lut_9_bit_4_fill;
wire [28:0] lut_9_bit_5_fill;
wire [28:0] lut_9_bit_6_fill;
wire [28:0] lut_9_bit_7_fill;
wire [28:0] lut_9_bit_8_fill;
wire [28:0] lut_9_bit_9_fill;
wire [28:0] lut_9_bit_10_fill;
wire [28:0] lut_9_bit_11_fill;
wire [28:0] lut_9_bit_12_fill;
wire [28:0] lut_9_bit_13_fill;
wire [28:0] lut_9_bit_14_fill;
wire [28:0] lut_9_bit_15_fill;
assign lut_9_bit_0_fill = {lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13], lut_val_9_n_0_pp[13],  lut_val_9_n_0_pp };
assign lut_9_bit_1_fill = {lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13], lut_val_9_n_1_pp[13],  lut_val_9_n_1_pp, 1'd0 };
assign lut_9_bit_2_fill = {lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13], lut_val_9_n_2_pp[13],  lut_val_9_n_2_pp, 2'd0 };
assign lut_9_bit_3_fill = {lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13], lut_val_9_n_3_pp[13],  lut_val_9_n_3_pp, 3'd0 };
assign lut_9_bit_4_fill = {lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13], lut_val_9_n_4_pp[13],  lut_val_9_n_4_pp, 4'd0 };
assign lut_9_bit_5_fill = {lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13], lut_val_9_n_5_pp[13],  lut_val_9_n_5_pp, 5'd0 };
assign lut_9_bit_6_fill = {lut_val_9_n_6_pp[13], lut_val_9_n_6_pp[13], lut_val_9_n_6_pp[13], lut_val_9_n_6_pp[13], lut_val_9_n_6_pp[13], lut_val_9_n_6_pp[13], lut_val_9_n_6_pp[13], lut_val_9_n_6_pp[13], lut_val_9_n_6_pp[13],  lut_val_9_n_6_pp, 6'd0 };
assign lut_9_bit_7_fill = {lut_val_9_n_7_pp[13], lut_val_9_n_7_pp[13], lut_val_9_n_7_pp[13], lut_val_9_n_7_pp[13], lut_val_9_n_7_pp[13], lut_val_9_n_7_pp[13], lut_val_9_n_7_pp[13], lut_val_9_n_7_pp[13],  lut_val_9_n_7_pp, 7'd0 };
assign lut_9_bit_8_fill = {lut_val_9_n_8_pp[13], lut_val_9_n_8_pp[13], lut_val_9_n_8_pp[13], lut_val_9_n_8_pp[13], lut_val_9_n_8_pp[13], lut_val_9_n_8_pp[13], lut_val_9_n_8_pp[13],  lut_val_9_n_8_pp, 8'd0 };
assign lut_9_bit_9_fill = {lut_val_9_n_9_pp[13], lut_val_9_n_9_pp[13], lut_val_9_n_9_pp[13], lut_val_9_n_9_pp[13], lut_val_9_n_9_pp[13], lut_val_9_n_9_pp[13],  lut_val_9_n_9_pp, 9'd0 };
assign lut_9_bit_10_fill = {lut_val_9_n_10_pp[13], lut_val_9_n_10_pp[13], lut_val_9_n_10_pp[13], lut_val_9_n_10_pp[13], lut_val_9_n_10_pp[13],  lut_val_9_n_10_pp, 10'd0 };
assign lut_9_bit_11_fill = {lut_val_9_n_11_pp[13], lut_val_9_n_11_pp[13], lut_val_9_n_11_pp[13], lut_val_9_n_11_pp[13],  lut_val_9_n_11_pp, 11'd0 };
assign lut_9_bit_12_fill = {lut_val_9_n_12_pp[13], lut_val_9_n_12_pp[13], lut_val_9_n_12_pp[13],  lut_val_9_n_12_pp, 12'd0 };
assign lut_9_bit_13_fill = {lut_val_9_n_13_pp[13], lut_val_9_n_13_pp[13],  lut_val_9_n_13_pp, 13'd0 };
assign lut_9_bit_14_fill = {lut_val_9_n_14_pp[13],  lut_val_9_n_14_pp, 14'd0 };
assign lut_9_bit_15_fill = { lut_val_9_n_15_pp, 15'd0 };
wire [29:0] tree_9_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_9_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_9_bit_0_fill), .bin(lut_9_bit_1_fill), .res(tree_9_pp_l_0_n_0_n) );
defparam Uadd_9_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_9_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_9_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_9_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_9_bit_2_fill), .bin(lut_9_bit_3_fill), .res(tree_9_pp_l_0_n_1_n) );
defparam Uadd_9_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_9_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_9_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_9_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_9_bit_4_fill), .bin(lut_9_bit_5_fill), .res(tree_9_pp_l_0_n_2_n) );
defparam Uadd_9_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_9_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_9_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_9_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_9_bit_6_fill), .bin(lut_9_bit_7_fill), .res(tree_9_pp_l_0_n_3_n) );
defparam Uadd_9_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_9_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_9_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_9_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_9_bit_8_fill), .bin(lut_9_bit_9_fill), .res(tree_9_pp_l_0_n_4_n) );
defparam Uadd_9_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_9_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_9_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_9_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_9_bit_10_fill), .bin(lut_9_bit_11_fill), .res(tree_9_pp_l_0_n_5_n) );
defparam Uadd_9_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_9_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_9_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_9_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_9_bit_12_fill), .bin(lut_9_bit_13_fill), .res(tree_9_pp_l_0_n_6_n) );
defparam Uadd_9_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_9_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_9_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_9_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_9_bit_14_fill), .bin(lut_9_bit_15_fill), .res(tree_9_pp_l_0_n_7_n) );
defparam Uadd_9_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_9_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_9_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_9_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_9_pp_l_0_n_0_n), .bin(tree_9_pp_l_0_n_1_n), .res(tree_9_pp_l_1_n_0_n) );
defparam Uadd_9_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_9_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_9_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_9_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_9_pp_l_0_n_2_n), .bin(tree_9_pp_l_0_n_3_n), .res(tree_9_pp_l_1_n_1_n) );
defparam Uadd_9_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_9_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_9_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_9_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_9_pp_l_0_n_4_n), .bin(tree_9_pp_l_0_n_5_n), .res(tree_9_pp_l_1_n_2_n) );
defparam Uadd_9_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_9_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_9_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_9_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_9_pp_l_0_n_6_n), .bin(tree_9_pp_l_0_n_7_n), .res(tree_9_pp_l_1_n_3_n) );
defparam Uadd_9_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_9_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_9_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_9_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_9_pp_l_1_n_0_n), .bin(tree_9_pp_l_1_n_1_n), .res(tree_9_pp_l_2_n_0_n) );
defparam Uadd_9_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_9_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_9_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_9_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_9_pp_l_1_n_2_n), .bin(tree_9_pp_l_1_n_3_n), .res(tree_9_pp_l_2_n_1_n) );
defparam Uadd_9_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_9_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_9_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_9_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_9_pp_l_2_n_0_n), .bin(tree_9_pp_l_2_n_1_n), .res(tree_9_pp_l_3_n_0_n) );
defparam Uadd_9_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_9_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_9_n;
assign lut_val_9_n=tree_9_pp_l_3_n_0_n;
wire [28:0] lut_10_bit_0_fill;
wire [28:0] lut_10_bit_1_fill;
wire [28:0] lut_10_bit_2_fill;
wire [28:0] lut_10_bit_3_fill;
wire [28:0] lut_10_bit_4_fill;
wire [28:0] lut_10_bit_5_fill;
wire [28:0] lut_10_bit_6_fill;
wire [28:0] lut_10_bit_7_fill;
wire [28:0] lut_10_bit_8_fill;
wire [28:0] lut_10_bit_9_fill;
wire [28:0] lut_10_bit_10_fill;
wire [28:0] lut_10_bit_11_fill;
wire [28:0] lut_10_bit_12_fill;
wire [28:0] lut_10_bit_13_fill;
wire [28:0] lut_10_bit_14_fill;
wire [28:0] lut_10_bit_15_fill;
assign lut_10_bit_0_fill = {lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13], lut_val_10_n_0_pp[13],  lut_val_10_n_0_pp };
assign lut_10_bit_1_fill = {lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13], lut_val_10_n_1_pp[13],  lut_val_10_n_1_pp, 1'd0 };
assign lut_10_bit_2_fill = {lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13], lut_val_10_n_2_pp[13],  lut_val_10_n_2_pp, 2'd0 };
assign lut_10_bit_3_fill = {lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13], lut_val_10_n_3_pp[13],  lut_val_10_n_3_pp, 3'd0 };
assign lut_10_bit_4_fill = {lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13], lut_val_10_n_4_pp[13],  lut_val_10_n_4_pp, 4'd0 };
assign lut_10_bit_5_fill = {lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13], lut_val_10_n_5_pp[13],  lut_val_10_n_5_pp, 5'd0 };
assign lut_10_bit_6_fill = {lut_val_10_n_6_pp[13], lut_val_10_n_6_pp[13], lut_val_10_n_6_pp[13], lut_val_10_n_6_pp[13], lut_val_10_n_6_pp[13], lut_val_10_n_6_pp[13], lut_val_10_n_6_pp[13], lut_val_10_n_6_pp[13], lut_val_10_n_6_pp[13],  lut_val_10_n_6_pp, 6'd0 };
assign lut_10_bit_7_fill = {lut_val_10_n_7_pp[13], lut_val_10_n_7_pp[13], lut_val_10_n_7_pp[13], lut_val_10_n_7_pp[13], lut_val_10_n_7_pp[13], lut_val_10_n_7_pp[13], lut_val_10_n_7_pp[13], lut_val_10_n_7_pp[13],  lut_val_10_n_7_pp, 7'd0 };
assign lut_10_bit_8_fill = {lut_val_10_n_8_pp[13], lut_val_10_n_8_pp[13], lut_val_10_n_8_pp[13], lut_val_10_n_8_pp[13], lut_val_10_n_8_pp[13], lut_val_10_n_8_pp[13], lut_val_10_n_8_pp[13],  lut_val_10_n_8_pp, 8'd0 };
assign lut_10_bit_9_fill = {lut_val_10_n_9_pp[13], lut_val_10_n_9_pp[13], lut_val_10_n_9_pp[13], lut_val_10_n_9_pp[13], lut_val_10_n_9_pp[13], lut_val_10_n_9_pp[13],  lut_val_10_n_9_pp, 9'd0 };
assign lut_10_bit_10_fill = {lut_val_10_n_10_pp[13], lut_val_10_n_10_pp[13], lut_val_10_n_10_pp[13], lut_val_10_n_10_pp[13], lut_val_10_n_10_pp[13],  lut_val_10_n_10_pp, 10'd0 };
assign lut_10_bit_11_fill = {lut_val_10_n_11_pp[13], lut_val_10_n_11_pp[13], lut_val_10_n_11_pp[13], lut_val_10_n_11_pp[13],  lut_val_10_n_11_pp, 11'd0 };
assign lut_10_bit_12_fill = {lut_val_10_n_12_pp[13], lut_val_10_n_12_pp[13], lut_val_10_n_12_pp[13],  lut_val_10_n_12_pp, 12'd0 };
assign lut_10_bit_13_fill = {lut_val_10_n_13_pp[13], lut_val_10_n_13_pp[13],  lut_val_10_n_13_pp, 13'd0 };
assign lut_10_bit_14_fill = {lut_val_10_n_14_pp[13],  lut_val_10_n_14_pp, 14'd0 };
assign lut_10_bit_15_fill = { lut_val_10_n_15_pp, 15'd0 };
wire [29:0] tree_10_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_10_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_10_bit_0_fill), .bin(lut_10_bit_1_fill), .res(tree_10_pp_l_0_n_0_n) );
defparam Uadd_10_lut_l_0_n_0_n.IN_WIDTH = 29;
defparam Uadd_10_lut_l_0_n_0_n.PIPE_DEPTH = 1;
wire [29:0] tree_10_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_10_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_10_bit_2_fill), .bin(lut_10_bit_3_fill), .res(tree_10_pp_l_0_n_1_n) );
defparam Uadd_10_lut_l_0_n_1_n.IN_WIDTH = 29;
defparam Uadd_10_lut_l_0_n_1_n.PIPE_DEPTH = 1;
wire [29:0] tree_10_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_10_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_10_bit_4_fill), .bin(lut_10_bit_5_fill), .res(tree_10_pp_l_0_n_2_n) );
defparam Uadd_10_lut_l_0_n_2_n.IN_WIDTH = 29;
defparam Uadd_10_lut_l_0_n_2_n.PIPE_DEPTH = 1;
wire [29:0] tree_10_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_10_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_10_bit_6_fill), .bin(lut_10_bit_7_fill), .res(tree_10_pp_l_0_n_3_n) );
defparam Uadd_10_lut_l_0_n_3_n.IN_WIDTH = 29;
defparam Uadd_10_lut_l_0_n_3_n.PIPE_DEPTH = 1;
wire [29:0] tree_10_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_10_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_10_bit_8_fill), .bin(lut_10_bit_9_fill), .res(tree_10_pp_l_0_n_4_n) );
defparam Uadd_10_lut_l_0_n_4_n.IN_WIDTH = 29;
defparam Uadd_10_lut_l_0_n_4_n.PIPE_DEPTH = 1;
wire [29:0] tree_10_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_10_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_10_bit_10_fill), .bin(lut_10_bit_11_fill), .res(tree_10_pp_l_0_n_5_n) );
defparam Uadd_10_lut_l_0_n_5_n.IN_WIDTH = 29;
defparam Uadd_10_lut_l_0_n_5_n.PIPE_DEPTH = 1;
wire [29:0] tree_10_pp_l_0_n_6_n;
sadd_lpm_cen Uadd_10_lut_l_0_n_6_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_10_bit_12_fill), .bin(lut_10_bit_13_fill), .res(tree_10_pp_l_0_n_6_n) );
defparam Uadd_10_lut_l_0_n_6_n.IN_WIDTH = 29;
defparam Uadd_10_lut_l_0_n_6_n.PIPE_DEPTH = 1;
wire [29:0] tree_10_pp_l_0_n_7_n;
sadd_lpm_cen Uadd_10_lut_l_0_n_7_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_10_bit_14_fill), .bin(lut_10_bit_15_fill), .res(tree_10_pp_l_0_n_7_n) );
defparam Uadd_10_lut_l_0_n_7_n.IN_WIDTH = 29;
defparam Uadd_10_lut_l_0_n_7_n.PIPE_DEPTH = 1;
wire [30:0] tree_10_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_10_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_10_pp_l_0_n_0_n), .bin(tree_10_pp_l_0_n_1_n), .res(tree_10_pp_l_1_n_0_n) );
defparam Uadd_10_lut_l_1_n_0_n.IN_WIDTH = 30;
defparam Uadd_10_lut_l_1_n_0_n.PIPE_DEPTH = 1;
wire [30:0] tree_10_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_10_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_10_pp_l_0_n_2_n), .bin(tree_10_pp_l_0_n_3_n), .res(tree_10_pp_l_1_n_1_n) );
defparam Uadd_10_lut_l_1_n_1_n.IN_WIDTH = 30;
defparam Uadd_10_lut_l_1_n_1_n.PIPE_DEPTH = 1;
wire [30:0] tree_10_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_10_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_10_pp_l_0_n_4_n), .bin(tree_10_pp_l_0_n_5_n), .res(tree_10_pp_l_1_n_2_n) );
defparam Uadd_10_lut_l_1_n_2_n.IN_WIDTH = 30;
defparam Uadd_10_lut_l_1_n_2_n.PIPE_DEPTH = 1;
wire [30:0] tree_10_pp_l_1_n_3_n;
sadd_lpm_cen Uadd_10_lut_l_1_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_10_pp_l_0_n_6_n), .bin(tree_10_pp_l_0_n_7_n), .res(tree_10_pp_l_1_n_3_n) );
defparam Uadd_10_lut_l_1_n_3_n.IN_WIDTH = 30;
defparam Uadd_10_lut_l_1_n_3_n.PIPE_DEPTH = 1;
wire [31:0] tree_10_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_10_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_10_pp_l_1_n_0_n), .bin(tree_10_pp_l_1_n_1_n), .res(tree_10_pp_l_2_n_0_n) );
defparam Uadd_10_lut_l_2_n_0_n.IN_WIDTH = 31;
defparam Uadd_10_lut_l_2_n_0_n.PIPE_DEPTH = 1;
wire [31:0] tree_10_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_10_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_10_pp_l_1_n_2_n), .bin(tree_10_pp_l_1_n_3_n), .res(tree_10_pp_l_2_n_1_n) );
defparam Uadd_10_lut_l_2_n_1_n.IN_WIDTH = 31;
defparam Uadd_10_lut_l_2_n_1_n.PIPE_DEPTH = 1;
wire [32:0] tree_10_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_10_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_10_pp_l_2_n_0_n), .bin(tree_10_pp_l_2_n_1_n), .res(tree_10_pp_l_3_n_0_n) );
defparam Uadd_10_lut_l_3_n_0_n.IN_WIDTH = 32;
defparam Uadd_10_lut_l_3_n_0_n.PIPE_DEPTH = 1;
wire [32:0] lut_val_10_n;
assign lut_val_10_n=tree_10_pp_l_3_n_0_n;
wire [33:0] fin_atree_l_0_n_0_n;
sadd_lpm_cen Uadd_cen_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_val_0_n), .bin(lut_val_1_n), .res(fin_atree_l_0_n_0_n) );
defparam Uadd_cen_l_0_n_0_n.IN_WIDTH = 33;
defparam Uadd_cen_l_0_n_0_n.PIPE_DEPTH = 1;
wire [33:0] fin_atree_l_0_n_1_n;
sadd_lpm_cen Uadd_cen_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_val_2_n), .bin(lut_val_3_n), .res(fin_atree_l_0_n_1_n) );
defparam Uadd_cen_l_0_n_1_n.IN_WIDTH = 33;
defparam Uadd_cen_l_0_n_1_n.PIPE_DEPTH = 1;
wire [33:0] fin_atree_l_0_n_2_n;
sadd_lpm_cen Uadd_cen_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_val_4_n), .bin(lut_val_5_n), .res(fin_atree_l_0_n_2_n) );
defparam Uadd_cen_l_0_n_2_n.IN_WIDTH = 33;
defparam Uadd_cen_l_0_n_2_n.PIPE_DEPTH = 1;
wire [33:0] fin_atree_l_0_n_3_n;
sadd_lpm_cen Uadd_cen_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_val_6_n), .bin(lut_val_7_n), .res(fin_atree_l_0_n_3_n) );
defparam Uadd_cen_l_0_n_3_n.IN_WIDTH = 33;
defparam Uadd_cen_l_0_n_3_n.PIPE_DEPTH = 1;
wire [33:0] fin_atree_l_0_n_4_n;
sadd_lpm_cen Uadd_cen_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_val_8_n), .bin(lut_val_9_n), .res(fin_atree_l_0_n_4_n) );
defparam Uadd_cen_l_0_n_4_n.IN_WIDTH = 33;
defparam Uadd_cen_l_0_n_4_n.PIPE_DEPTH = 1;
wire [33:0] fin_atree_l_0_n_5_n;
sadd_lpm_cen Uadd_cen_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_val_10_n), .bin(33'd0), .res(fin_atree_l_0_n_5_n) );
defparam Uadd_cen_l_0_n_5_n.IN_WIDTH = 33;
defparam Uadd_cen_l_0_n_5_n.PIPE_DEPTH = 1;
wire [34:0] fin_atree_l_1_n_0_n;
sadd_lpm_cen Uadd_cen_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(fin_atree_l_0_n_0_n), .bin(fin_atree_l_0_n_1_n), .res(fin_atree_l_1_n_0_n) );
defparam Uadd_cen_l_1_n_0_n.IN_WIDTH = 34;
defparam Uadd_cen_l_1_n_0_n.PIPE_DEPTH = 1;
wire [34:0] fin_atree_l_1_n_1_n;
sadd_lpm_cen Uadd_cen_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(fin_atree_l_0_n_2_n), .bin(fin_atree_l_0_n_3_n), .res(fin_atree_l_1_n_1_n) );
defparam Uadd_cen_l_1_n_1_n.IN_WIDTH = 34;
defparam Uadd_cen_l_1_n_1_n.PIPE_DEPTH = 1;
wire [34:0] fin_atree_l_1_n_2_n;
sadd_lpm_cen Uadd_cen_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(fin_atree_l_0_n_4_n), .bin(fin_atree_l_0_n_5_n), .res(fin_atree_l_1_n_2_n) );
defparam Uadd_cen_l_1_n_2_n.IN_WIDTH = 34;
defparam Uadd_cen_l_1_n_2_n.PIPE_DEPTH = 1;
wire [35:0] fin_atree_l_2_n_0_n;
sadd_lpm_cen Uadd_cen_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(fin_atree_l_1_n_0_n), .bin(fin_atree_l_1_n_1_n), .res(fin_atree_l_2_n_0_n) );
defparam Uadd_cen_l_2_n_0_n.IN_WIDTH = 35;
defparam Uadd_cen_l_2_n_0_n.PIPE_DEPTH = 1;
wire [35:0] fin_atree_l_2_n_1_n;
sadd_lpm_cen Uadd_cen_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(fin_atree_l_1_n_2_n), .bin(35'd0), .res(fin_atree_l_2_n_1_n) );
defparam Uadd_cen_l_2_n_1_n.IN_WIDTH = 35;
defparam Uadd_cen_l_2_n_1_n.PIPE_DEPTH = 1;
wire [36:0] fin_atree_l_3_n_0_n;
sadd_lpm_cen Uadd_cen_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(fin_atree_l_2_n_0_n), .bin(fin_atree_l_2_n_1_n), .res(fin_atree_l_3_n_0_n) );
defparam Uadd_cen_l_3_n_0_n.IN_WIDTH = 36;
defparam Uadd_cen_l_3_n_0_n.PIPE_DEPTH = 1;
wire [36:0] mac_res;
assign mac_res=fin_atree_l_3_n_0_n;
wire [36:0] atree_res;
mac_tl Umtl (.clk(clk),
             .data_in(mac_res),
             .data_out(atree_res));
defparam Umtl.DATA_WIDTH = 37;
wire [30:0] fir_int_res;
assign fir_int_res = atree_res [30:0];
wire [30:0]fir_int_res_fill;
assign fir_int_res_fill =  fir_int_res[30 :0];
parameter TOT_WIDTH = ACCUM_WIDTH;
assign fir_result = fir_int_res_fill[TOT_WIDTH-MSB_RM-1:LSB_RM];
wire pre_rdy;
assign rdy_to_ld = pre_rdy;
assign done = done_int;
par_ctrl Uctrl(.rst(rst),
		.clk(clk),
		.clk_en(clk_en),
		.done(done_int),
		.rdy_int(rdy_int),
		.rdy_to_ld(pre_rdy));
defparam Uctrl.REG_LEN = 11;
defparam Uctrl.REG_BIT = 4;
defparam Uctrl.CH_WIDTH =0;
defparam Uctrl.NUM_CH =1;
endmodule