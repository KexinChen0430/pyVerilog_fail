module simulation done. ***");
      $finish;
    end // aes_core_test
endmodule