module OUTBUF (
	input D,
	(* iopad_external_pin *)
	output PAD
);
	assign PAD = D;
endmodule