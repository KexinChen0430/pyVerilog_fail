module arrayed_wire;
   wire [3:0][7:0] n2;
endmodule