module bug868 (ifmp);
   if_bug777.master ifmp;
endmodule