module b14 (
  clock,
  reset,
  addr,
  datai,
  datao,
  rd,
  wr
)
;
input clock ;
input reset ;
output [19:0] addr ;
input [31:0] datai ;
output [31:0] datao ;
output rd ;
output wr ;
wire clock ;
wire reset ;
wire rd ;
wire wr ;
wire [0:0] state;
wire [31:0] ir;
wire [28:0] reg3;
wire [31:0] ir_3;
wire [31:0] reg2;
wire [31:0] m_2;
wire [31:0] reg1;
wire [31:0] r_4;
wire [31:0] reg0;
wire [30:0] un11_r_cry;
wire [1:0] d;
wire [30:30] r_6;
wire [30:0] un26_r_cry;
wire [31:0] reg2_16;
wire [19:0] un1_inf_abs0_10;
wire [19:0] un1_inf_abs0_11;
wire [18:0] reg0_28;
wire [18:0] reg1_16;
wire [28:0] reg3_17;
wire [28:0] b18_cry;
wire [30:30] r_4_3_lut6_2_O5;
wire [9:0] un14_r_0_data_tmp;
wire [16:1] t_6;
wire [0:0] d_cnst;
wire [0:0] dce;
wire [31:0] inf_abs0_2;
wire [31:1] reg3_1_1;
wire [31:0] t_1;
wire [18:17] reg0_28_7_a1;
wire [24:24] reg0_28_7_d;
wire [24:21] reg3_17_a0;
wire [29:29] reg2_16_11_a1;
wire [29:17] reg2_16_11_a2;
wire [29:17] reg2_16_11_a3;
wire [1:0] r_4_2_a0;
wire [13:13] reg3_17_4_a2;
wire [10:10] r_4_1_RNIDBOH1;
wire [25:21] reg2_16_11_a4;
wire [9:9] r_4_1_RNIS3K91;
wire [7:7] r_4_1_RNIFO731;
wire [8:8] r_4_1_RNIIQ731;
wire [5:5] r_4_1_RNI9K731;
wire [6:6] r_4_1_RNICM731;
wire [3:3] r_4_2_a1_lut6_2_RNI5V8R3;
wire [3:3] r_4_2_a1_lut6_2_RNI2T8R3;
wire [24:21] \d_cnst_sn.reg3_17_0_tz ;
wire [4:0] \d_cnst_sn.r_4_0_0 ;
wire [20:20] reg2_16_2_d;
wire [3:3] r_4_2_a1_lut6_2_O6;
wire [3:3] r_4_2_a1_lut6_2_O5;
wire [28:28] \d_cnst_sn.reg2_16_0_1_tz ;
wire [28:28] \d_cnst_sn.reg2_16_11_1_tz ;
wire [7:7] \d_cnst_sn.reg0_28_a0_1 ;
wire [5:5] \d_cnst_sn.reg1_16_a2_0 ;
wire [4:4] \d_cnst_sn.reg0_28_a1_1 ;
wire [3:3] \d_cnst_sn.reg1_16_a0_1 ;
wire [9:9] \d_cnst_sn.reg0_28_7_a0_0 ;
wire [24:24] \d_cnst_sn.reg3_17_a1_2 ;
wire [0:0] state_i;
wire [31:31] r_4_i;
wire [31:0] m_2_i;
wire [28:20] \d_cnst_sn.reg3_17_4_a2_0 ;
wire [21:21] \d_cnst_sn.reg3_17_a2_2_0 ;
wire [8:2] \d_cnst_sn.reg0_1 ;
wire [8:3] \d_cnst_sn.reg1_1 ;
wire [28:12] \d_cnst_sn.reg3_17_6_0 ;
wire [19:12] \d_cnst_sn.reg3_17_6_1 ;
wire [20:19] \d_cnst_sn.reg0_28_0 ;
wire [25:20] \d_cnst_sn.reg2_16_0 ;
wire [29:20] \d_cnst_sn.reg2_16_1 ;
wire [17:17] \d_cnst_sn.reg0_0 ;
wire [18:18] \d_cnst_sn.reg1_0 ;
wire [28:26] \d_cnst_sn.reg2_16_0_1_0 ;
wire [31:31] r_4_3_ci;
wire [31:31] ir_fast;
wire [31:31] ir_3_fast;
wire [31:31] inf_abs0_2_0;
wire [31:31] inf_abs0_2_1;
wire [1:1] \d_cnst_sn.reg2_16_11muxnet_0 ;
wire [1:1] \d_cnst_sn.reg2_16_11muxnet_1 ;
wire b ;
wire VCC ;
wire GND ;
wire addr_4_sqmuxa_1 ;
wire un14_r_0_I_83 ;
wire b18 ;
wire un11_reg0_s_1 ;
wire un11_reg0_s_2 ;
wire un11_reg0_s_3 ;
wire un11_reg0_s_4 ;
wire un11_reg0_s_5 ;
wire un11_reg0_s_6 ;
wire un11_reg0_s_7 ;
wire un11_reg0_s_8 ;
wire un11_reg0_s_9 ;
wire un11_reg0_s_10 ;
wire un11_reg0_s_11 ;
wire un11_reg0_s_12 ;
wire un11_reg0_s_13 ;
wire un11_reg0_s_14 ;
wire un11_reg0_s_15 ;
wire un11_reg0_s_16 ;
wire un11_reg0_s_17 ;
wire un11_reg0_s_18 ;
wire un11_reg0_s_19 ;
wire un11_reg0_s_20 ;
wire un11_reg0_s_21 ;
wire un11_reg0_s_22 ;
wire un11_reg0_s_23 ;
wire un11_reg0_s_24 ;
wire un11_reg0_s_25 ;
wire un11_reg0_s_26 ;
wire un11_reg0_s_27 ;
wire un11_reg0_s_28 ;
wire un11_reg0_s_29 ;
wire rd_18 ;
wire un11_r_df0 ;
wire un11_r_lt0 ;
wire un11_r_df2 ;
wire un11_r_lt2 ;
wire un11_r_df4 ;
wire un11_r_lt4 ;
wire un11_r_df6 ;
wire un11_r_lt6 ;
wire un11_r_df8 ;
wire un11_r_lt8 ;
wire un11_r_df10 ;
wire un11_r_lt10 ;
wire un11_r_df12 ;
wire un11_r_lt12 ;
wire un11_r_df14 ;
wire un11_r_lt14 ;
wire un11_r_df16 ;
wire un11_r_lt16 ;
wire un11_r_df18 ;
wire un11_r_lt18 ;
wire un11_r_df20 ;
wire un11_r_lt20 ;
wire un11_r_df22 ;
wire un11_r_lt22 ;
wire un11_r_df24 ;
wire un11_r_lt24 ;
wire un11_r_df26 ;
wire un11_r_lt26 ;
wire un11_r_df28 ;
wire un11_r_lt28 ;
wire un11_r_df30 ;
wire un11_r_lt30 ;
wire b18_df0 ;
wire b18_lt0 ;
wire b18_df2 ;
wire b18_lt2 ;
wire b18_df4 ;
wire b18_lt4 ;
wire b18_df6 ;
wire b18_lt6 ;
wire b18_df8 ;
wire b18_lt8 ;
wire b18_df10 ;
wire b18_lt10 ;
wire b18_df12 ;
wire b18_lt12 ;
wire b18_df14 ;
wire b18_lt14 ;
wire b18_df16 ;
wire b18_lt16 ;
wire b18_df18 ;
wire b18_lt18 ;
wire b18_df20 ;
wire b18_lt20 ;
wire b18_df22 ;
wire b18_lt22 ;
wire b18_df24 ;
wire b18_lt24 ;
wire b18_df26 ;
wire b18_lt26 ;
wire b18_df28 ;
wire b18_lt28 ;
wire b18_df30 ;
wire b18_lt30 ;
wire un26_r_df0 ;
wire un26_r_lt0 ;
wire un26_r_df2 ;
wire un26_r_lt2 ;
wire un26_r_df4 ;
wire un26_r_lt4 ;
wire un26_r_df6 ;
wire un26_r_lt6 ;
wire un26_r_df8 ;
wire un26_r_lt8 ;
wire un26_r_df10 ;
wire un26_r_lt10 ;
wire un26_r_df12 ;
wire un26_r_lt12 ;
wire un26_r_df14 ;
wire un26_r_lt14 ;
wire un26_r_df16 ;
wire un26_r_lt16 ;
wire un26_r_df18 ;
wire un26_r_lt18 ;
wire un26_r_df20 ;
wire un26_r_lt20 ;
wire un26_r_df22 ;
wire un26_r_lt22 ;
wire un26_r_df24 ;
wire un26_r_lt24 ;
wire un26_r_df26 ;
wire un26_r_lt26 ;
wire un26_r_df28 ;
wire un26_r_lt28 ;
wire un26_r_df30 ;
wire un26_r_lt30 ;
wire r_4_3_30_680_i_m2 ;
wire r_4_3_29_706_i_m2 ;
wire r_4_3_28_732_i_m2 ;
wire r_4_3_27_758_i_m2 ;
wire r_4_3_25_810_i_m2 ;
wire r_4_3_24_836_i_m2 ;
wire r_4_3_23_1078_i_m2 ;
wire r_4_3_22_1104_i_m2 ;
wire r_4_3_20_1156_i_m2 ;
wire r_4_3_19_1182_i_m2 ;
wire r_4_3_18_1208_i_m2 ;
wire r_4_3_17_1234_i_m2 ;
wire r_4_3_16_1260_i_m2 ;
wire r_4_3_15_1286_i_m2 ;
wire r_4_3_14_1312_i_m2 ;
wire r_4_3_13_1338_i_m2 ;
wire r_4_3_12_1364_i_m2 ;
wire r_4_3_11_1390_i_m2 ;
wire r_4_3_10_1416_i_m2 ;
wire r_4_3_9_1442_i_m2 ;
wire r_4_3_8_1467 ;
wire r_4_3_6_1508_i_m2 ;
wire r_4_3_5_1534_i_m2 ;
wire r_4_3_4_1560_i_m2 ;
wire r_4_3_3_1586_i_m2 ;
wire r_4_3_2_1612_i_m2 ;
wire r_4_3_1_1638_i_m2 ;
wire r_4_3_0_1664_i_m2 ;
wire r_4_3_1690_i_m2 ;
wire reg1_16_9 ;
wire reg1_16_8_1837 ;
wire reg1_16_7_1870 ;
wire reg0_28_10_2261_a6_3_2_lut6_2_RNIOK9O5 ;
wire reg0_28_8_2327 ;
wire reg0_28_7_2360 ;
wire reg0_28_6_2393 ;
wire reg0_28_5_2426 ;
wire reg0_28_4_2459 ;
wire reg0_28_3_2492 ;
wire un14_r_0_N_2 ;
wire un14_r_0_N_7 ;
wire un14_r_0_N_14 ;
wire un14_r_0_N_21 ;
wire un14_r_0_N_28 ;
wire un14_r_0_N_35 ;
wire un14_r_0_N_42 ;
wire un14_r_0_N_49 ;
wire un14_r_0_N_56 ;
wire un14_r_0_N_63 ;
wire un14_r_0_N_70 ;
wire N_28 ;
wire N_3550 ;
wire N_3856 ;
wire N_2724 ;
wire N_3673 ;
wire N_939 ;
wire N_3_0 ;
wire N_971 ;
wire N_13 ;
wire un1_cf ;
wire N_1688 ;
wire reg3_1_sqmuxa ;
wire un1_df_16 ;
wire N_1750 ;
wire reg3_14_sqmuxa ;
wire N_1812 ;
wire N_1810 ;
wire N_1841 ;
wire N_1661 ;
wire N_1816 ;
wire N_1681 ;
wire N_1743 ;
wire N_938 ;
wire N_970 ;
wire N_1033 ;
wire N_513_i ;
wire N_3873_2 ;
wire N_512_i ;
wire un1_df_1 ;
wire un36_df ;
wire d_cnst_sm0 ;
wire N_3913 ;
wire N_1342 ;
wire N_1374 ;
wire N_514_i ;
wire N_1566 ;
wire N_1584 ;
wire N_1890 ;
wire un86_df ;
wire N_1664 ;
wire N_1819 ;
wire N_1682 ;
wire N_1837 ;
wire N_527_i ;
wire N_1042 ;
wire N_3916 ;
wire N_1270 ;
wire N_1132 ;
wire N_1892 ;
wire N_2641 ;
wire un87_df ;
wire N_7_i ;
wire N_1043 ;
wire b_2_sqmuxa ;
wire N_3912 ;
wire N_895 ;
wire N_526_i ;
wire un1_df_17_2 ;
wire N_1493 ;
wire N_1337 ;
wire N_1343 ;
wire N_1369 ;
wire N_1375 ;
wire N_1561 ;
wire N_1567 ;
wire N_934 ;
wire N_2722 ;
wire N_45 ;
wire N_54 ;
wire m7 ;
wire N_1901 ;
wire addr_4_sqmuxa_1_1 ;
wire un1_b57 ;
wire rd_4_sqmuxa ;
wire N_1740 ;
wire N_2240_i ;
wire N_3568 ;
wire N_2660_2 ;
wire N_915 ;
wire N_919 ;
wire N_918 ;
wire N_1076 ;
wire N_1044 ;
wire N_953 ;
wire N_921 ;
wire N_959 ;
wire N_927 ;
wire N_969 ;
wire N_937 ;
wire N_1084 ;
wire N_1052 ;
wire N_965 ;
wire N_933 ;
wire N_1741 ;
wire N_1679 ;
wire N_1742 ;
wire N_1680 ;
wire N_3614 ;
wire N_974 ;
wire N_942 ;
wire N_1838 ;
wire N_1683 ;
wire N_1039 ;
wire N_1085 ;
wire N_1053 ;
wire N_1083 ;
wire N_1051 ;
wire N_1040 ;
wire N_1038 ;
wire N_952 ;
wire N_920 ;
wire N_1077 ;
wire N_1045 ;
wire N_1081 ;
wire N_1049 ;
wire N_1827 ;
wire N_1672 ;
wire N_1082 ;
wire N_1050 ;
wire N_964 ;
wire N_932 ;
wire N_962 ;
wire N_930 ;
wire N_967 ;
wire N_935 ;
wire N_1079 ;
wire N_1047 ;
wire N_1068 ;
wire N_1036 ;
wire N_1078 ;
wire N_1046 ;
wire N_968 ;
wire N_936 ;
wire N_1069 ;
wire N_1037 ;
wire N_916 ;
wire N_1080 ;
wire N_1048 ;
wire N_1815 ;
wire N_1660 ;
wire N_1820 ;
wire N_1818 ;
wire N_1814 ;
wire N_1665 ;
wire N_1663 ;
wire N_1659 ;
wire N_1752 ;
wire N_1690 ;
wire N_955 ;
wire N_923 ;
wire N_954 ;
wire N_922 ;
wire N_1823 ;
wire N_1668 ;
wire N_956 ;
wire N_924 ;
wire N_1822 ;
wire N_1667 ;
wire N_957 ;
wire N_925 ;
wire N_1829 ;
wire N_1824 ;
wire N_1674 ;
wire N_1669 ;
wire N_961 ;
wire N_929 ;
wire N_1817 ;
wire N_1662 ;
wire N_963 ;
wire N_931 ;
wire N_1830 ;
wire N_1826 ;
wire N_1675 ;
wire N_1671 ;
wire N_960 ;
wire N_928 ;
wire N_1832 ;
wire N_1677 ;
wire N_1831 ;
wire N_1821 ;
wire N_1676 ;
wire N_1666 ;
wire N_1041 ;
wire N_1828 ;
wire N_1673 ;
wire N_972 ;
wire N_940 ;
wire N_1840 ;
wire N_1685 ;
wire N_975 ;
wire N_943 ;
wire N_1839 ;
wire N_1684 ;
wire N_973 ;
wire N_941 ;
wire N_958 ;
wire N_926 ;
wire un1_b59 ;
wire N_1813 ;
wire N_1732 ;
wire N_1670 ;
wire N_1658 ;
wire N_1751 ;
wire N_1689 ;
wire N_1583 ;
wire N_1582 ;
wire N_1581 ;
wire N_1580 ;
wire N_1575 ;
wire N_1574 ;
wire N_1573 ;
wire N_1572 ;
wire N_1571 ;
wire N_1570 ;
wire N_1569 ;
wire N_1568 ;
wire N_1565 ;
wire N_1564 ;
wire N_1563 ;
wire N_1562 ;
wire N_1560 ;
wire N_1035 ;
wire N_1363 ;
wire N_1362 ;
wire N_1361 ;
wire N_1354 ;
wire N_1353 ;
wire N_1352 ;
wire N_1351 ;
wire N_1383 ;
wire N_1350 ;
wire N_1382 ;
wire N_1349 ;
wire N_1381 ;
wire N_1348 ;
wire N_1380 ;
wire N_1347 ;
wire N_1379 ;
wire N_1346 ;
wire N_1378 ;
wire N_1345 ;
wire N_1377 ;
wire N_1344 ;
wire N_1376 ;
wire N_1341 ;
wire N_1373 ;
wire N_1340 ;
wire N_1372 ;
wire N_1339 ;
wire N_1371 ;
wire N_1338 ;
wire N_1370 ;
wire N_1336 ;
wire N_1368 ;
wire N_1335 ;
wire inf_abs0_2_axb_0 ;
wire inf_abs0_2_cry_0 ;
wire inf_abs0_2_axb_1 ;
wire inf_abs0_2_cry_1 ;
wire inf_abs0_2_axb_2 ;
wire inf_abs0_2_cry_2 ;
wire inf_abs0_2_axb_3 ;
wire inf_abs0_2_cry_3 ;
wire inf_abs0_2_axb_4 ;
wire inf_abs0_2_cry_4 ;
wire inf_abs0_2_axb_5 ;
wire inf_abs0_2_cry_5 ;
wire inf_abs0_2_axb_6 ;
wire inf_abs0_2_cry_6 ;
wire inf_abs0_2_axb_7 ;
wire inf_abs0_2_cry_7 ;
wire inf_abs0_2_axb_8 ;
wire inf_abs0_2_cry_8 ;
wire inf_abs0_2_axb_9 ;
wire inf_abs0_2_cry_9 ;
wire inf_abs0_2_axb_10 ;
wire inf_abs0_2_cry_10 ;
wire inf_abs0_2_axb_11 ;
wire inf_abs0_2_cry_11 ;
wire inf_abs0_2_axb_12 ;
wire inf_abs0_2_cry_12 ;
wire inf_abs0_2_axb_13 ;
wire inf_abs0_2_cry_13 ;
wire inf_abs0_2_axb_14 ;
wire inf_abs0_2_cry_14 ;
wire inf_abs0_2_axb_15 ;
wire inf_abs0_2_cry_15 ;
wire inf_abs0_2_axb_16 ;
wire inf_abs0_2_cry_16 ;
wire inf_abs0_2_axb_17 ;
wire inf_abs0_2_cry_17 ;
wire inf_abs0_2_axb_18 ;
wire inf_abs0_2_cry_18 ;
wire inf_abs0_2_axb_19 ;
wire inf_abs0_2_cry_19 ;
wire inf_abs0_2_axb_20 ;
wire inf_abs0_2_cry_20 ;
wire inf_abs0_2_axb_21 ;
wire inf_abs0_2_cry_21 ;
wire inf_abs0_2_axb_22 ;
wire inf_abs0_2_cry_22 ;
wire inf_abs0_2_axb_23 ;
wire inf_abs0_2_cry_23 ;
wire inf_abs0_2_axb_24 ;
wire inf_abs0_2_cry_24 ;
wire inf_abs0_2_axb_25 ;
wire inf_abs0_2_cry_25 ;
wire inf_abs0_2_axb_26 ;
wire inf_abs0_2_cry_26 ;
wire inf_abs0_2_axb_27 ;
wire inf_abs0_2_cry_27 ;
wire inf_abs0_2_axb_28 ;
wire inf_abs0_2_cry_28 ;
wire inf_abs0_2_axb_29 ;
wire inf_abs0_2_cry_29 ;
wire inf_abs0_2_axb_30 ;
wire reg3_1_1_axb_0 ;
wire reg3_1_1_cry_0 ;
wire reg3_1_1_axb_1 ;
wire reg3_1_1_cry_1 ;
wire reg3_1_1_axb_2 ;
wire reg3_1_1_cry_2 ;
wire reg3_1_1_axb_3 ;
wire reg3_1_1_cry_3 ;
wire reg3_1_1_axb_4 ;
wire reg3_1_1_cry_4 ;
wire reg3_1_1_axb_5 ;
wire reg3_1_1_cry_5 ;
wire reg3_1_1_axb_6 ;
wire reg3_1_1_cry_6 ;
wire reg3_1_1_axb_7 ;
wire reg3_1_1_cry_7 ;
wire reg3_1_1_axb_8 ;
wire reg3_1_1_cry_8 ;
wire reg3_1_1_axb_9 ;
wire reg3_1_1_cry_9 ;
wire reg3_1_1_axb_10 ;
wire reg3_1_1_cry_10 ;
wire reg3_1_1_axb_11 ;
wire reg3_1_1_cry_11 ;
wire reg3_1_1_axb_12 ;
wire reg3_1_1_cry_12 ;
wire reg3_1_1_axb_13 ;
wire reg3_1_1_cry_13 ;
wire reg3_1_1_axb_14 ;
wire reg3_1_1_cry_14 ;
wire reg3_1_1_axb_15 ;
wire reg3_1_1_cry_15 ;
wire reg3_1_1_axb_16 ;
wire reg3_1_1_cry_16 ;
wire reg3_1_1_axb_17 ;
wire reg3_1_1_cry_17 ;
wire reg3_1_1_axb_18 ;
wire reg3_1_1_cry_18 ;
wire reg3_1_1_axb_19 ;
wire reg3_1_1_cry_19 ;
wire reg3_1_1_cry_20 ;
wire reg3_1_1_cry_21 ;
wire reg3_1_1_cry_22 ;
wire reg3_1_1_cry_23 ;
wire reg3_1_1_cry_24 ;
wire reg3_1_1_cry_25 ;
wire reg3_1_1_cry_26 ;
wire reg3_1_1_cry_27 ;
wire reg3_1_1_cry_28 ;
wire reg3_1_1_axb_29 ;
wire reg3_1_1_cry_29 ;
wire reg3_1_1_axb_30 ;
wire reg3_1_1_cry_30 ;
wire reg3_1_1_axb_31 ;
wire un3_t_s_1 ;
wire un3_t_s_2 ;
wire un3_t_s_3 ;
wire un3_t_s_4 ;
wire un3_t_s_5 ;
wire un3_t_s_6 ;
wire un3_t_s_7 ;
wire un3_t_s_8 ;
wire un3_t_s_9 ;
wire un3_t_s_10 ;
wire un3_t_s_11 ;
wire un3_t_s_12 ;
wire un3_t_s_13 ;
wire un3_t_s_14 ;
wire un3_t_s_15 ;
wire un3_t_s_16 ;
wire un3_t_s_17 ;
wire un3_t_s_18 ;
wire un3_t_s_19 ;
wire un3_t_s_20 ;
wire un3_t_s_21 ;
wire un3_t_s_22 ;
wire un3_t_s_23 ;
wire un3_t_s_24 ;
wire un3_t_s_25 ;
wire un3_t_s_26 ;
wire un3_t_s_27 ;
wire un3_t_s_28 ;
wire un3_t_s_29 ;
wire un3_t_s_30 ;
wire un3_t_s_31 ;
wire un3_t_cry_0 ;
wire un3_t_cry_1 ;
wire un3_t_axb_2 ;
wire un3_t_cry_2 ;
wire un3_t_cry_3 ;
wire un3_t_cry_4 ;
wire un3_t_cry_5 ;
wire un3_t_cry_6 ;
wire un3_t_cry_7 ;
wire un3_t_cry_8 ;
wire un3_t_cry_9 ;
wire un3_t_cry_10 ;
wire un3_t_cry_11 ;
wire un3_t_cry_12 ;
wire un3_t_cry_13 ;
wire un3_t_cry_14 ;
wire un3_t_cry_15 ;
wire un3_t_cry_16 ;
wire un3_t_cry_17 ;
wire un3_t_cry_18 ;
wire un3_t_cry_19 ;
wire un3_t_cry_20 ;
wire un3_t_cry_21 ;
wire un3_t_cry_22 ;
wire un3_t_cry_23 ;
wire un3_t_cry_24 ;
wire un3_t_cry_25 ;
wire un3_t_cry_26 ;
wire un3_t_cry_27 ;
wire un3_t_cry_28 ;
wire un3_t_axb_29 ;
wire un3_t_cry_29 ;
wire un3_t_axb_30 ;
wire un3_t_cry_30 ;
wire un3_t_axb_31 ;
wire un11_reg0_axb_0 ;
wire un11_reg0_cry_0 ;
wire un11_reg0_axb_1 ;
wire un11_reg0_cry_1 ;
wire un11_reg0_axb_2 ;
wire un11_reg0_cry_2 ;
wire un11_reg0_axb_3 ;
wire un11_reg0_cry_3 ;
wire un11_reg0_axb_4 ;
wire un11_reg0_cry_4 ;
wire un11_reg0_axb_5 ;
wire un11_reg0_cry_5 ;
wire un11_reg0_axb_6 ;
wire un11_reg0_cry_6 ;
wire un11_reg0_axb_7 ;
wire un11_reg0_cry_7 ;
wire un11_reg0_axb_8 ;
wire un11_reg0_cry_8 ;
wire un11_reg0_axb_9 ;
wire un11_reg0_cry_9 ;
wire un11_reg0_axb_10 ;
wire un11_reg0_cry_10 ;
wire un11_reg0_axb_11 ;
wire un11_reg0_cry_11 ;
wire un11_reg0_axb_12 ;
wire un11_reg0_cry_12 ;
wire un11_reg0_axb_13 ;
wire un11_reg0_cry_13 ;
wire un11_reg0_axb_14 ;
wire un11_reg0_cry_14 ;
wire un11_reg0_axb_15 ;
wire un11_reg0_cry_15 ;
wire un11_reg0_axb_16 ;
wire un11_reg0_cry_16 ;
wire un11_reg0_axb_17 ;
wire un11_reg0_cry_17 ;
wire un11_reg0_axb_18 ;
wire un11_reg0_cry_18 ;
wire un11_reg0_axb_19 ;
wire un11_reg0_cry_19 ;
wire un11_reg0_axb_20 ;
wire un11_reg0_cry_20 ;
wire un11_reg0_axb_21 ;
wire un11_reg0_cry_21 ;
wire un11_reg0_axb_22 ;
wire un11_reg0_cry_22 ;
wire un11_reg0_axb_23 ;
wire un11_reg0_cry_23 ;
wire un11_reg0_axb_24 ;
wire un11_reg0_cry_24 ;
wire un11_reg0_axb_25 ;
wire un11_reg0_cry_25 ;
wire un11_reg0_axb_26 ;
wire un11_reg0_cry_26 ;
wire un11_reg0_axb_27 ;
wire un11_reg0_cry_27 ;
wire un11_reg0_axb_28 ;
wire un11_reg0_cry_28 ;
wire un11_reg0_axb_29 ;
wire un32_reg0_s_1 ;
wire un32_reg0_s_2 ;
wire un32_reg0_s_3 ;
wire un32_reg0_s_4 ;
wire un32_reg0_s_5 ;
wire un32_reg0_s_6 ;
wire un32_reg0_s_7 ;
wire un32_reg0_s_8 ;
wire un32_reg0_s_9 ;
wire un32_reg0_s_10 ;
wire un32_reg0_s_11 ;
wire un32_reg0_s_12 ;
wire un32_reg0_s_13 ;
wire un32_reg0_s_14 ;
wire un32_reg0_s_15 ;
wire un32_reg0_s_16 ;
wire un32_reg0_s_17 ;
wire un32_reg0_s_18 ;
wire un32_reg0_s_19 ;
wire un32_reg0_s_20 ;
wire un32_reg0_s_21 ;
wire un32_reg0_s_22 ;
wire un32_reg0_s_23 ;
wire un32_reg0_s_24 ;
wire un32_reg0_s_25 ;
wire un32_reg0_s_26 ;
wire un32_reg0_s_27 ;
wire un32_reg0_s_28 ;
wire un32_reg0_s_29 ;
wire un32_reg0_cry_0 ;
wire un32_reg0_axb_1 ;
wire un32_reg0_cry_1 ;
wire un32_reg0_axb_2 ;
wire un32_reg0_cry_2 ;
wire un32_reg0_axb_3 ;
wire un32_reg0_cry_3 ;
wire un32_reg0_axb_4 ;
wire un32_reg0_cry_4 ;
wire un32_reg0_axb_5 ;
wire un32_reg0_cry_5 ;
wire un32_reg0_axb_6 ;
wire un32_reg0_cry_6 ;
wire un32_reg0_axb_7 ;
wire un32_reg0_cry_7 ;
wire un32_reg0_axb_8 ;
wire un32_reg0_cry_8 ;
wire un32_reg0_axb_9 ;
wire un32_reg0_cry_9 ;
wire un32_reg0_axb_10 ;
wire un32_reg0_cry_10 ;
wire un32_reg0_axb_11 ;
wire un32_reg0_cry_11 ;
wire un32_reg0_axb_12 ;
wire un32_reg0_cry_12 ;
wire un32_reg0_axb_13 ;
wire un32_reg0_cry_13 ;
wire un32_reg0_axb_14 ;
wire un32_reg0_cry_14 ;
wire un32_reg0_axb_15 ;
wire un32_reg0_cry_15 ;
wire un32_reg0_axb_16 ;
wire un32_reg0_cry_16 ;
wire un32_reg0_axb_17 ;
wire un32_reg0_cry_17 ;
wire un32_reg0_axb_18 ;
wire un32_reg0_cry_18 ;
wire un32_reg0_axb_19 ;
wire un32_reg0_cry_19 ;
wire un32_reg0_axb_20 ;
wire un32_reg0_cry_20 ;
wire un32_reg0_axb_21 ;
wire un32_reg0_cry_21 ;
wire un32_reg0_axb_22 ;
wire un32_reg0_cry_22 ;
wire un32_reg0_axb_23 ;
wire un32_reg0_cry_23 ;
wire un32_reg0_axb_24 ;
wire un32_reg0_cry_24 ;
wire un32_reg0_axb_25 ;
wire un32_reg0_cry_25 ;
wire un32_reg0_axb_26 ;
wire un32_reg0_cry_26 ;
wire un32_reg0_axb_27 ;
wire un32_reg0_cry_27 ;
wire un32_reg0_axb_28 ;
wire un32_reg0_cry_28 ;
wire un32_reg0_axb_29 ;
wire un1_inf_abs0_cry_0 ;
wire un1_inf_abs0_axb_1 ;
wire un1_inf_abs0_cry_1 ;
wire un1_inf_abs0_axb_2 ;
wire un1_inf_abs0_cry_2 ;
wire un1_inf_abs0_axb_3 ;
wire un1_inf_abs0_cry_3 ;
wire un1_inf_abs0_axb_4 ;
wire un1_inf_abs0_cry_4 ;
wire un1_inf_abs0_axb_5 ;
wire un1_inf_abs0_cry_5 ;
wire un1_inf_abs0_axb_6 ;
wire un1_inf_abs0_cry_6 ;
wire un1_inf_abs0_axb_7 ;
wire un1_inf_abs0_cry_7 ;
wire un1_inf_abs0_axb_8 ;
wire un1_inf_abs0_cry_8 ;
wire un1_inf_abs0_axb_9 ;
wire un1_inf_abs0_cry_9 ;
wire un1_inf_abs0_axb_10 ;
wire un1_inf_abs0_cry_10 ;
wire un1_inf_abs0_axb_11 ;
wire un1_inf_abs0_cry_11 ;
wire un1_inf_abs0_axb_12 ;
wire un1_inf_abs0_cry_12 ;
wire un1_inf_abs0_axb_13 ;
wire un1_inf_abs0_cry_13 ;
wire un1_inf_abs0_axb_14 ;
wire un1_inf_abs0_cry_14 ;
wire un1_inf_abs0_axb_15 ;
wire un1_inf_abs0_cry_15 ;
wire un1_inf_abs0_axb_16 ;
wire un1_inf_abs0_cry_16 ;
wire un1_inf_abs0_axb_17 ;
wire un1_inf_abs0_cry_17 ;
wire un1_inf_abs0_axb_18 ;
wire un1_inf_abs0_cry_18 ;
wire un1_inf_abs0_axb_19 ;
wire un1_inf_abs0_0_cry_0 ;
wire un1_inf_abs0_0_axb_1 ;
wire un1_inf_abs0_0_cry_1 ;
wire un1_inf_abs0_0_axb_2 ;
wire un1_inf_abs0_0_cry_2 ;
wire un1_inf_abs0_0_axb_3 ;
wire un1_inf_abs0_0_cry_3 ;
wire un1_inf_abs0_0_axb_4 ;
wire un1_inf_abs0_0_cry_4 ;
wire un1_inf_abs0_0_axb_5 ;
wire un1_inf_abs0_0_cry_5 ;
wire un1_inf_abs0_0_axb_6 ;
wire un1_inf_abs0_0_cry_6 ;
wire un1_inf_abs0_0_axb_7 ;
wire un1_inf_abs0_0_cry_7 ;
wire un1_inf_abs0_0_axb_8 ;
wire un1_inf_abs0_0_cry_8 ;
wire un1_inf_abs0_0_axb_9 ;
wire un1_inf_abs0_0_cry_9 ;
wire un1_inf_abs0_0_axb_10 ;
wire un1_inf_abs0_0_cry_10 ;
wire un1_inf_abs0_0_axb_11 ;
wire un1_inf_abs0_0_cry_11 ;
wire un1_inf_abs0_0_axb_12 ;
wire un1_inf_abs0_0_cry_12 ;
wire un1_inf_abs0_0_axb_13 ;
wire un1_inf_abs0_0_cry_13 ;
wire un1_inf_abs0_0_axb_14 ;
wire un1_inf_abs0_0_cry_14 ;
wire un1_inf_abs0_0_axb_15 ;
wire un1_inf_abs0_0_cry_15 ;
wire un1_inf_abs0_0_axb_16 ;
wire un1_inf_abs0_0_cry_16 ;
wire un1_inf_abs0_0_axb_17 ;
wire un1_inf_abs0_0_cry_17 ;
wire un1_inf_abs0_0_axb_18 ;
wire un1_inf_abs0_0_cry_18 ;
wire un1_inf_abs0_0_axb_19 ;
wire un3_reg3_s_1 ;
wire un3_reg3_s_2 ;
wire un3_reg3_s_3 ;
wire un3_reg3_s_4 ;
wire un3_reg3_s_5 ;
wire un3_reg3_s_6 ;
wire un3_reg3_s_7 ;
wire un3_reg3_s_8 ;
wire un3_reg3_s_9 ;
wire un3_reg3_s_10 ;
wire un3_reg3_s_11 ;
wire un3_reg3_s_12 ;
wire un3_reg3_s_13 ;
wire un3_reg3_s_14 ;
wire un3_reg3_s_15 ;
wire un3_reg3_s_16 ;
wire un3_reg3_s_17 ;
wire un3_reg3_s_18 ;
wire un3_reg3_s_19 ;
wire un3_reg3_s_20 ;
wire un3_reg3_s_21 ;
wire un3_reg3_s_22 ;
wire un3_reg3_s_23 ;
wire un3_reg3_s_24 ;
wire un3_reg3_s_25 ;
wire un3_reg3_cry_25 ;
wire un3_reg3_axb_1 ;
wire un3_reg3_cry_1 ;
wire un3_reg3_axb_2 ;
wire un3_reg3_cry_2 ;
wire un3_reg3_axb_3 ;
wire un3_reg3_cry_3 ;
wire un3_reg3_axb_4 ;
wire un3_reg3_cry_4 ;
wire un3_reg3_axb_5 ;
wire un3_reg3_cry_5 ;
wire un3_reg3_axb_6 ;
wire un3_reg3_cry_6 ;
wire un3_reg3_axb_7 ;
wire un3_reg3_cry_7 ;
wire un3_reg3_axb_8 ;
wire un3_reg3_cry_8 ;
wire un3_reg3_axb_9 ;
wire un3_reg3_cry_9 ;
wire un3_reg3_axb_10 ;
wire un3_reg3_cry_10 ;
wire un3_reg3_axb_11 ;
wire un3_reg3_cry_11 ;
wire un3_reg3_axb_12 ;
wire un3_reg3_cry_12 ;
wire un3_reg3_axb_13 ;
wire un3_reg3_cry_13 ;
wire un3_reg3_axb_14 ;
wire un3_reg3_cry_14 ;
wire un3_reg3_axb_15 ;
wire un3_reg3_cry_15 ;
wire un3_reg3_axb_16 ;
wire un3_reg3_cry_16 ;
wire un3_reg3_axb_17 ;
wire un3_reg3_cry_17 ;
wire un3_reg3_axb_18 ;
wire un3_reg3_cry_18 ;
wire un3_reg3_axb_19 ;
wire un3_reg3_cry_19 ;
wire un3_reg3_axb_20 ;
wire un3_reg3_cry_20 ;
wire un3_reg3_axb_21 ;
wire un3_reg3_cry_21 ;
wire un3_reg3_axb_22 ;
wire un3_reg3_cry_22 ;
wire un3_reg3_axb_23 ;
wire un3_reg3_cry_23 ;
wire un3_reg3_axb_24 ;
wire un3_reg3_cry_24 ;
wire un3_reg3_axb_25 ;
wire t_1_cry_0 ;
wire t_1_cry_1 ;
wire t_1_cry_2 ;
wire t_1_cry_3 ;
wire t_1_cry_4 ;
wire t_1_cry_5 ;
wire t_1_cry_6 ;
wire t_1_cry_7 ;
wire t_1_cry_8 ;
wire t_1_cry_9 ;
wire t_1_cry_10 ;
wire t_1_cry_11 ;
wire t_1_cry_12 ;
wire t_1_cry_13 ;
wire t_1_cry_14 ;
wire t_1_cry_15 ;
wire t_1_cry_16 ;
wire t_1_cry_17 ;
wire t_1_cry_18 ;
wire t_1_cry_19 ;
wire t_1_cry_20 ;
wire t_1_cry_21 ;
wire t_1_cry_22 ;
wire t_1_cry_23 ;
wire t_1_cry_24 ;
wire t_1_cry_25 ;
wire t_1_cry_26 ;
wire t_1_cry_27 ;
wire t_1_cry_28 ;
wire t_1_cry_29 ;
wire t_1_cry_30 ;
wire \d_cnst_sn.reg1_16_8_1837_2_tz  ;
wire reg0_28_sn_m6_lut6_2_O5 ;
wire \d_cnst_sn.reg3_17_sn_m7_0  ;
wire reg3_1_sqmuxa_RNIH1DM1 ;
wire reg3_1_sqmuxa_RNIE1DM1 ;
wire reg3_1_sqmuxa_RNIQMUH1 ;
wire reg3_1_sqmuxa_RNITMUH1 ;
wire reg3_1_sqmuxa_RNIKMUH1 ;
wire reg3_1_sqmuxa_RNINMUH1 ;
wire reg3_1_sqmuxa_RNIHMUH1 ;
wire reg3_1_sqmuxa_RNIEMUH1 ;
wire reg0_m9_i_a1 ;
wire \d_cnst_sn.reg2_N_3_mux  ;
wire g0_2_0_i2_lut6_2_O6 ;
wire reg3_N_7_i_RNO ;
wire \d_cnst_sn.reg1_16_9_1804_3_tz  ;
wire \d_cnst_sn.addr_20_iv_1052_i_a6_1_0  ;
wire \d_cnst_sn.reg0_m8_e_0  ;
wire \d_cnst_sn.reg3_5_sqmuxa_2_1  ;
wire \d_cnst_sn.reg0_28_9_2294_a6_3_0  ;
wire N_3910 ;
wire \d_cnst_sn.un1_state_3_1  ;
wire \d_cnst_sn.b60_0  ;
wire \d_cnst_sn.b64_0  ;
wire \d_cnst_sn.reg0_m9_i_a3_0  ;
wire reg3_17_sn_N_5 ;
wire \d_cnst_sn.reg0_28_2526_a5_1_0  ;
wire N_4571_i ;
wire N_4570_i ;
wire N_4569_i ;
wire N_4568_i ;
wire N_4567_i ;
wire N_4566_i ;
wire N_4565_i ;
wire N_4564_i ;
wire N_4563_i ;
wire N_4562_i ;
wire N_4561_i ;
wire N_4560_i ;
wire N_4559_i ;
wire N_4558_i ;
wire N_4557_i ;
wire N_4556_i ;
wire N_4555_i ;
wire N_4554_i ;
wire N_4553_i ;
wire N_4552_i ;
wire N_4551_i ;
wire N_4550_i ;
wire N_4549_i ;
wire N_4548_i ;
wire N_4547_i ;
wire N_4546_i ;
wire N_4545_i ;
wire N_4544_i ;
wire N_4543_i ;
wire N_4542_i ;
wire N_4541_i ;
wire \d_cnst_sn.reg3_N_7_i  ;
wire N_2099_i ;
wire addr_0_sqmuxa_1_i ;
wire N_2119_i ;
wire N_2139_i ;
wire N_2159_i ;
wire N_2179_i ;
wire N_2199_i ;
wire N_2219_i ;
wire N_56_i ;
wire N_2267_i ;
wire N_47_i ;
wire N_2315_i ;
wire N_2335_i ;
wire N_36_i ;
wire N_2516_i ;
wire N_2536_i ;
wire N_2556_i ;
wire N_2576_i ;
wire N_2596_i ;
wire N_2616_i ;
wire N_2636_i ;
wire N_2656_i ;
wire un1_state_1_0_i ;
wire un1_state_3_i ;
wire un1_state_4_i ;
wire \d_cnst_sn.addr_20_iv_1052_i_a6_2_0  ;
wire \d_cnst_sn.m26_0_1  ;
wire \d_cnst_sn.m19_0_1  ;
wire \d_cnst_sn.addr_20_iv_7_654_i_1  ;
wire \d_cnst_sn.addr_20_iv_8_627_i_1  ;
wire \d_cnst_sn.addr_20_iv_16_389_i_1  ;
wire \d_cnst_sn.addr_20_iv_12_497_i_1  ;
wire \d_cnst_sn.addr_20_iv_10_562_i_1  ;
wire \d_cnst_sn.addr_20_iv_14_443_i_2  ;
wire \d_cnst_sn.addr_20_iv_15_416_i_1  ;
wire \d_cnst_sn.addr_20_iv_17_362_i_1  ;
wire \d_cnst_sn.addr_20_iv_13_470_i_1  ;
wire \d_cnst_sn.addr_20_iv_18_335_i_1  ;
wire \d_cnst_sn.addr_20_iv_2_971_i_0  ;
wire \d_cnst_sn.addr_20_iv_1_998_i_0  ;
wire \d_cnst_sn.addr_20_iv_1052_i_0  ;
wire \d_cnst_sn.addr_20_iv_0_1025_i_0  ;
wire \d_cnst_sn.addr_20_iv_3_944_i_0  ;
wire \d_cnst_sn.addr_20_iv_4_917_i_0  ;
wire \d_cnst_sn.addr_20_iv_5_890_i_0  ;
wire \d_cnst_sn.addr_20_iv_6_863_i_0  ;
wire \d_cnst_sn.reg0_28_12_2195_a6_1_2_0  ;
wire \d_cnst_sn.reg0_m9_i_a0_0  ;
wire \d_cnst_sn.reg0_28_5_2426_a6_1_1  ;
wire \d_cnst_sn.reg0_28_5_2426_3_1  ;
wire \d_cnst_sn.reg0_28_8_2327_a6_1_1  ;
wire \d_cnst_sn.reg0_28_6_2393_3_1  ;
wire \d_cnst_sn.reg0_28_6_2393_a6_1_1  ;
wire \d_cnst_sn.reg0_28_7_2360_3_1  ;
wire \d_cnst_sn.reg0_28_7_2360_a6_1_1  ;
wire \d_cnst_sn.reg0_28_14_2135_1_a0_2  ;
wire \d_cnst_sn.reg0_28_9_2294_a6_1_1  ;
wire \d_cnst_sn.reg0_28_9_2294_3_1  ;
wire \d_cnst_sn.reg1_16_7_1870_3_1  ;
wire \d_cnst_sn.reg0_28_10_2261_a6_1_1  ;
wire \d_cnst_sn.reg1_16_8_1837_3_1  ;
wire \d_cnst_sn.reg0_28_11_2228_a6_1_1  ;
wire \d_cnst_sn.reg0_28_3_2492_0  ;
wire \d_cnst_sn.reg0_28_3_2492_1  ;
wire \d_cnst_sn.reg0_28_4_2459_0  ;
wire \d_cnst_sn.reg0_28_8_2327_0  ;
wire \d_cnst_sn.reg0_28_5_2426_0  ;
wire \d_cnst_sn.reg0_28_6_2393_0  ;
wire \d_cnst_sn.reg0_28_7_2360_0  ;
wire \d_cnst_sn.reg0_28_14_0  ;
wire \d_cnst_sn.reg0_28_9_2294_0  ;
wire \d_cnst_sn.reg1_16_7_1870_0  ;
wire \d_cnst_sn.reg1_16_8_1837_0  ;
wire b_0 ;
wire un3_t_axb_28 ;
wire un3_t_axb_27 ;
wire un3_t_axb_26 ;
wire un3_t_axb_25 ;
wire un3_t_axb_24 ;
wire un3_t_axb_23 ;
wire un3_t_axb_22 ;
wire un3_t_axb_21 ;
wire un3_t_axb_20 ;
wire un3_t_axb_19 ;
wire un3_t_axb_18 ;
wire un3_t_axb_17 ;
wire un3_t_axb_16 ;
wire un3_t_axb_15 ;
wire un3_t_axb_14 ;
wire un3_t_axb_13 ;
wire un3_t_axb_12 ;
wire un3_t_axb_11 ;
wire un3_t_axb_10 ;
wire un3_t_axb_9 ;
wire un3_t_axb_8 ;
wire un3_t_axb_7 ;
wire un3_t_axb_6 ;
wire un3_t_axb_5 ;
wire un3_t_axb_4 ;
wire un3_t_axb_3 ;
wire un3_t_axb_1 ;
wire un3_t_axb_0 ;
wire reg3_1_1_axb_28 ;
wire reg3_1_1_axb_27 ;
wire reg3_1_1_axb_26 ;
wire reg3_1_1_axb_25 ;
wire reg3_1_1_axb_24 ;
wire reg3_1_1_axb_23 ;
wire reg3_1_1_axb_22 ;
wire reg3_1_1_axb_21 ;
wire reg3_1_1_axb_20 ;
wire t_1_cry_0_cy ;
wire un3_t_cry_0_cy ;
wire N_7 ;
wire N_12 ;
wire \d_cnst_sn.g0_3_a2_2  ;
wire \d_cnst_sn.g0_3_1  ;
wire \d_cnst_sn.g3  ;
wire \d_cnst_sn.reg0_N_13_0  ;
wire \d_cnst_sn.g0_0_2  ;
wire \d_cnst_sn.g0_1  ;
wire N_7_0 ;
wire \d_cnst_sn.g0_0_0_a5_0_0  ;
wire \d_cnst_sn.g0_0_0_a5_2  ;
wire \d_cnst_sn.g0_0_0_1  ;
wire N_3856_rep1 ;
wire N_3569_rep1 ;
wire N_3289_rep1 ;
wire N_3315_rep1 ;
wire N_3550_rep1 ;
wire N_3341_rep1 ;
wire N_3673_rep1 ;
wire N_3699_rep1 ;
wire N_3725_rep1 ;
wire N_3751_rep1 ;
wire N_3777_rep1 ;
wire N_3803_rep1 ;
wire N_3829_rep1 ;
wire \d_cnst_sn.g0_rn_1  ;
wire reg0_28_7_rep1 ;
wire d_cnst_ss0_x ;
wire un1_cf_x ;
wire un3_reg3_cry_25_0 ;
wire un3_reg3_cry_25_1 ;
wire inf_abs0_2_cry_29_0 ;
wire inf_abs0_2_cry_29_1 ;
  GND GND_cZ (
	.G(GND)
);
  VCC VCC_cZ (
	.P(VCC)
);
// @7:74
  MUXF8 \d_cnst_sn.reg2_16_11mux[1]  (
	.I0(\d_cnst_sn.reg2_16_11muxnet_0 [1]),
	.I1(\d_cnst_sn.reg2_16_11muxnet_1 [1]),
	.S(N_513_i),
	.O(reg2_16[1])
);
  MUXF7 \d_cnst_sn.reg2_16_11mux_RNO_0[1]  (
	.I0(N_1560),
	.I1(t_6[1]),
	.S(N_514_i),
	.O(\d_cnst_sn.reg2_16_11muxnet_1 [1])
);
  MUXF7 \d_cnst_sn.reg2_16_11mux_RNO[1]  (
	.I0(N_1336),
	.I1(N_1368),
	.S(N_514_i),
	.O(\d_cnst_sn.reg2_16_11muxnet_0 [1])
);
// @7:83
  LUT1 inf_abs0_2_cry_29_outextlut (
	.I0(VCC),
	.O(inf_abs0_2_cry_29_1)
);
defparam inf_abs0_2_cry_29_outextlut.INIT=2'h3;
// @7:95
  LUT1 un3_reg3_cry_25_outextlut (
	.I0(VCC),
	.O(un3_reg3_cry_25_1)
);
defparam un3_reg3_cry_25_outextlut.INIT=2'h3;
// @7:83
  LUT1 inf_abs0_2_cry_30_outextlut (
	.I0(VCC),
	.O(inf_abs0_2_1[31])
);
defparam inf_abs0_2_cry_30_outextlut.INIT=2'h3;
// @7:97
  LUT6_2 \d_cnst_sn.r_4_3_lut6_2[30]  (
	.I0(reg0[30]),
	.I1(reg1[30]),
	.I2(reg2[30]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(inf_abs0_2[31]),
	.O6(r_4[30]),
	.O5(r_4_3_lut6_2_O5[30])
);
defparam \d_cnst_sn.r_4_3_lut6_2[30] .INIT=64'hAAAAAAAA00F0CCAA;
// @7:118
  LUT4 un11_r_df0_cZ (
	.I0(m_2[0]),
	.I1(m_2[1]),
	.I2(r_4[0]),
	.I3(r_4[1]),
	.O(un11_r_df0)
);
defparam un11_r_df0_cZ.INIT=16'h8421;
// @7:118
  LUT4 un11_r_df2_cZ (
	.I0(N_28),
	.I1(m_2[2]),
	.I2(m_2[3]),
	.I3(r_4[3]),
	.O(un11_r_df2)
);
defparam un11_r_df2_cZ.INIT=16'h9009;
// @7:118
  LUT4 un11_r_df4_cZ (
	.I0(m_2[4]),
	.I1(m_2[5]),
	.I2(r_4[4]),
	.I3(r_4[5]),
	.O(un11_r_df4)
);
defparam un11_r_df4_cZ.INIT=16'h8421;
// @7:118
  LUT4 un11_r_df6_cZ (
	.I0(m_2[6]),
	.I1(m_2[7]),
	.I2(r_4[6]),
	.I3(r_4[7]),
	.O(un11_r_df6)
);
defparam un11_r_df6_cZ.INIT=16'h8421;
// @7:118
  LUT4 un11_r_df8_cZ (
	.I0(m_2[8]),
	.I1(m_2[9]),
	.I2(r_4[8]),
	.I3(r_4[9]),
	.O(un11_r_df8)
);
defparam un11_r_df8_cZ.INIT=16'h8421;
// @7:118
  LUT4 un11_r_df10_cZ (
	.I0(m_2[10]),
	.I1(m_2[11]),
	.I2(r_4[10]),
	.I3(r_4[11]),
	.O(un11_r_df10)
);
defparam un11_r_df10_cZ.INIT=16'h8421;
// @7:118
  LUT4 un11_r_df12_cZ (
	.I0(m_2[12]),
	.I1(m_2[13]),
	.I2(r_4[12]),
	.I3(r_4[13]),
	.O(un11_r_df12)
);
defparam un11_r_df12_cZ.INIT=16'h8421;
// @7:118
  LUT4 un11_r_df14_cZ (
	.I0(m_2[14]),
	.I1(m_2[15]),
	.I2(r_4[14]),
	.I3(r_4[15]),
	.O(un11_r_df14)
);
defparam un11_r_df14_cZ.INIT=16'h8421;
// @7:118
  LUT4 un11_r_df16_cZ (
	.I0(m_2[16]),
	.I1(m_2[17]),
	.I2(r_4[16]),
	.I3(r_4[17]),
	.O(un11_r_df16)
);
defparam un11_r_df16_cZ.INIT=16'h8421;
// @7:118
  LUT4 un11_r_df18_cZ (
	.I0(m_2[18]),
	.I1(m_2[19]),
	.I2(r_4[18]),
	.I3(r_4[19]),
	.O(un11_r_df18)
);
defparam un11_r_df18_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df0_cZ (
	.I0(m_2[0]),
	.I1(m_2[1]),
	.I2(r_4[0]),
	.I3(r_4[1]),
	.O(b18_df0)
);
defparam b18_df0_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df2_cZ (
	.I0(N_28),
	.I1(m_2[2]),
	.I2(m_2[3]),
	.I3(r_4[3]),
	.O(b18_df2)
);
defparam b18_df2_cZ.INIT=16'h9009;
// @7:143
  LUT4 b18_df4_cZ (
	.I0(m_2[4]),
	.I1(m_2[5]),
	.I2(r_4[4]),
	.I3(r_4[5]),
	.O(b18_df4)
);
defparam b18_df4_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df6_cZ (
	.I0(m_2[6]),
	.I1(m_2[7]),
	.I2(r_4[6]),
	.I3(r_4[7]),
	.O(b18_df6)
);
defparam b18_df6_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df8_cZ (
	.I0(m_2[8]),
	.I1(m_2[9]),
	.I2(r_4[8]),
	.I3(r_4[9]),
	.O(b18_df8)
);
defparam b18_df8_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df10_cZ (
	.I0(m_2[10]),
	.I1(m_2[11]),
	.I2(r_4[10]),
	.I3(r_4[11]),
	.O(b18_df10)
);
defparam b18_df10_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df12_cZ (
	.I0(m_2[12]),
	.I1(m_2[13]),
	.I2(r_4[12]),
	.I3(r_4[13]),
	.O(b18_df12)
);
defparam b18_df12_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df14_cZ (
	.I0(m_2[14]),
	.I1(m_2[15]),
	.I2(r_4[14]),
	.I3(r_4[15]),
	.O(b18_df14)
);
defparam b18_df14_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df16_cZ (
	.I0(m_2[16]),
	.I1(m_2[17]),
	.I2(r_4[16]),
	.I3(r_4[17]),
	.O(b18_df16)
);
defparam b18_df16_cZ.INIT=16'h8421;
// @7:143
  LUT4 b18_df18_cZ (
	.I0(m_2[18]),
	.I1(m_2[19]),
	.I2(r_4[18]),
	.I3(r_4[19]),
	.O(b18_df18)
);
defparam b18_df18_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df0_cZ (
	.I0(m_2[0]),
	.I1(m_2[1]),
	.I2(r_4[0]),
	.I3(r_4[1]),
	.O(un26_r_df0)
);
defparam un26_r_df0_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df2_cZ (
	.I0(N_28),
	.I1(m_2[2]),
	.I2(m_2[3]),
	.I3(r_4[3]),
	.O(un26_r_df2)
);
defparam un26_r_df2_cZ.INIT=16'h9009;
// @7:151
  LUT4 un26_r_df4_cZ (
	.I0(m_2[4]),
	.I1(m_2[5]),
	.I2(r_4[4]),
	.I3(r_4[5]),
	.O(un26_r_df4)
);
defparam un26_r_df4_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df6_cZ (
	.I0(m_2[6]),
	.I1(m_2[7]),
	.I2(r_4[6]),
	.I3(r_4[7]),
	.O(un26_r_df6)
);
defparam un26_r_df6_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df8_cZ (
	.I0(m_2[8]),
	.I1(m_2[9]),
	.I2(r_4[8]),
	.I3(r_4[9]),
	.O(un26_r_df8)
);
defparam un26_r_df8_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df10_cZ (
	.I0(m_2[10]),
	.I1(m_2[11]),
	.I2(r_4[10]),
	.I3(r_4[11]),
	.O(un26_r_df10)
);
defparam un26_r_df10_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df12_cZ (
	.I0(m_2[12]),
	.I1(m_2[13]),
	.I2(r_4[12]),
	.I3(r_4[13]),
	.O(un26_r_df12)
);
defparam un26_r_df12_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df14_cZ (
	.I0(m_2[14]),
	.I1(m_2[15]),
	.I2(r_4[14]),
	.I3(r_4[15]),
	.O(un26_r_df14)
);
defparam un26_r_df14_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df16_cZ (
	.I0(m_2[16]),
	.I1(m_2[17]),
	.I2(r_4[16]),
	.I3(r_4[17]),
	.O(un26_r_df16)
);
defparam un26_r_df16_cZ.INIT=16'h8421;
// @7:151
  LUT4 un26_r_df18_cZ (
	.I0(m_2[18]),
	.I1(m_2[19]),
	.I2(r_4[18]),
	.I3(r_4[19]),
	.O(un26_r_df18)
);
defparam un26_r_df18_cZ.INIT=16'h8421;
// @7:83
  LUT2 inf_abs0_2_axb_0_cZ (
	.I0(ir[0]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_0)
);
defparam inf_abs0_2_axb_0_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_1_cZ (
	.I0(ir[1]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_1)
);
defparam inf_abs0_2_axb_1_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_2_cZ (
	.I0(ir[2]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_2)
);
defparam inf_abs0_2_axb_2_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_3_cZ (
	.I0(ir[3]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_3)
);
defparam inf_abs0_2_axb_3_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_4_cZ (
	.I0(ir[4]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_4)
);
defparam inf_abs0_2_axb_4_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_5_cZ (
	.I0(ir[5]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_5)
);
defparam inf_abs0_2_axb_5_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_6_cZ (
	.I0(ir[6]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_6)
);
defparam inf_abs0_2_axb_6_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_7_cZ (
	.I0(ir[7]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_7)
);
defparam inf_abs0_2_axb_7_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_8_cZ (
	.I0(ir[8]),
	.I1(ir_fast[31]),
	.O(inf_abs0_2_axb_8)
);
defparam inf_abs0_2_axb_8_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_9_cZ (
	.I0(ir[9]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_9)
);
defparam inf_abs0_2_axb_9_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_10_cZ (
	.I0(ir[10]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_10)
);
defparam inf_abs0_2_axb_10_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_11_cZ (
	.I0(ir[11]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_11)
);
defparam inf_abs0_2_axb_11_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_12_cZ (
	.I0(ir[12]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_12)
);
defparam inf_abs0_2_axb_12_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_13_cZ (
	.I0(ir[13]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_13)
);
defparam inf_abs0_2_axb_13_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_14_cZ (
	.I0(ir[14]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_14)
);
defparam inf_abs0_2_axb_14_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_15_cZ (
	.I0(ir[15]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_15)
);
defparam inf_abs0_2_axb_15_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_16_cZ (
	.I0(ir[16]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_16)
);
defparam inf_abs0_2_axb_16_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_17_cZ (
	.I0(ir[17]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_17)
);
defparam inf_abs0_2_axb_17_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_18_cZ (
	.I0(ir[18]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_18)
);
defparam inf_abs0_2_axb_18_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_19_cZ (
	.I0(ir[19]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_19)
);
defparam inf_abs0_2_axb_19_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_20_cZ (
	.I0(ir[20]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_20)
);
defparam inf_abs0_2_axb_20_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_21_cZ (
	.I0(ir[21]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_21)
);
defparam inf_abs0_2_axb_21_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_22_cZ (
	.I0(ir[22]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_22)
);
defparam inf_abs0_2_axb_22_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_23_cZ (
	.I0(ir[23]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_23)
);
defparam inf_abs0_2_axb_23_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_24_cZ (
	.I0(ir[24]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_24)
);
defparam inf_abs0_2_axb_24_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_25_cZ (
	.I0(ir[25]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_25)
);
defparam inf_abs0_2_axb_25_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_26_cZ (
	.I0(ir[26]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_26)
);
defparam inf_abs0_2_axb_26_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_27_cZ (
	.I0(ir[27]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_27)
);
defparam inf_abs0_2_axb_27_cZ.INIT=4'h6;
// @7:83
  LUT2 inf_abs0_2_axb_28_cZ (
	.I0(ir[28]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_28)
);
defparam inf_abs0_2_axb_28_cZ.INIT=4'h6;
  LUT4 \datai_RNI2UAU[20]  (
	.I0(datai[20]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_20)
);
defparam \datai_RNI2UAU[20] .INIT=16'hFF57;
  LUT4 \datai_RNI3VAU[21]  (
	.I0(datai[21]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_21)
);
defparam \datai_RNI3VAU[21] .INIT=16'hFF57;
  LUT4 \datai_RNI40BU[22]  (
	.I0(datai[22]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_22)
);
defparam \datai_RNI40BU[22] .INIT=16'hFF57;
  LUT4 \datai_RNI51BU[23]  (
	.I0(datai[23]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_23)
);
defparam \datai_RNI51BU[23] .INIT=16'hFF57;
  LUT4 \datai_RNI62BU[24]  (
	.I0(datai[24]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_24)
);
defparam \datai_RNI62BU[24] .INIT=16'hFF57;
  LUT4 \datai_RNI73BU[25]  (
	.I0(datai[25]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_25)
);
defparam \datai_RNI73BU[25] .INIT=16'hFF57;
  LUT4 \datai_RNI84BU[26]  (
	.I0(datai[26]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_26)
);
defparam \datai_RNI84BU[26] .INIT=16'hFF57;
  LUT4 \datai_RNI95BU[27]  (
	.I0(datai[27]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_27)
);
defparam \datai_RNI95BU[27] .INIT=16'hFF57;
  LUT4 \datai_RNIA6BU[28]  (
	.I0(datai[28]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_28)
);
defparam \datai_RNIA6BU[28] .INIT=16'hFF57;
// @7:243
  LUT4 reg3_1_1_axb_29_cZ (
	.I0(datai[29]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_29)
);
defparam reg3_1_1_axb_29_cZ.INIT=16'hFF57;
// @7:243
  LUT4 reg3_1_1_axb_30_cZ (
	.I0(datai[30]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[31]),
	.O(reg3_1_1_axb_30)
);
defparam reg3_1_1_axb_30_cZ.INIT=16'hFF57;
// @7:74
  LUT2 un1_inf_abs0_cry_0_RNO (
	.I0(inf_abs0_2[0]),
	.I1(reg2[0]),
	.O(un1_inf_abs0_10[0])
);
defparam un1_inf_abs0_cry_0_RNO.INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIEGHO[1]  (
	.I0(inf_abs0_2[1]),
	.I1(reg2[1]),
	.O(un1_inf_abs0_axb_1)
);
defparam \reg2_RNIEGHO[1] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIGHHO[2]  (
	.I0(inf_abs0_2[2]),
	.I1(reg2[2]),
	.O(un1_inf_abs0_axb_2)
);
defparam \reg2_RNIGHHO[2] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIIIHO[3]  (
	.I0(inf_abs0_2[3]),
	.I1(reg2[3]),
	.O(un1_inf_abs0_axb_3)
);
defparam \reg2_RNIIIHO[3] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIKJHO[4]  (
	.I0(inf_abs0_2[4]),
	.I1(reg2[4]),
	.O(un1_inf_abs0_axb_4)
);
defparam \reg2_RNIKJHO[4] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIMKHO[5]  (
	.I0(inf_abs0_2[5]),
	.I1(reg2[5]),
	.O(un1_inf_abs0_axb_5)
);
defparam \reg2_RNIMKHO[5] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIOLHO[6]  (
	.I0(inf_abs0_2[6]),
	.I1(reg2[6]),
	.O(un1_inf_abs0_axb_6)
);
defparam \reg2_RNIOLHO[6] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIQMHO[7]  (
	.I0(inf_abs0_2[7]),
	.I1(reg2[7]),
	.O(un1_inf_abs0_axb_7)
);
defparam \reg2_RNIQMHO[7] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNISNHO[8]  (
	.I0(inf_abs0_2[8]),
	.I1(reg2[8]),
	.O(un1_inf_abs0_axb_8)
);
defparam \reg2_RNISNHO[8] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIUOHO[9]  (
	.I0(inf_abs0_2[9]),
	.I1(reg2[9]),
	.O(un1_inf_abs0_axb_9)
);
defparam \reg2_RNIUOHO[9] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIEK0A[10]  (
	.I0(inf_abs0_2[10]),
	.I1(reg2[10]),
	.O(un1_inf_abs0_axb_10)
);
defparam \reg2_RNIEK0A[10] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIGL0A[11]  (
	.I0(inf_abs0_2[11]),
	.I1(reg2[11]),
	.O(un1_inf_abs0_axb_11)
);
defparam \reg2_RNIGL0A[11] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIIM0A[12]  (
	.I0(inf_abs0_2[12]),
	.I1(reg2[12]),
	.O(un1_inf_abs0_axb_12)
);
defparam \reg2_RNIIM0A[12] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIKN0A[13]  (
	.I0(inf_abs0_2[13]),
	.I1(reg2[13]),
	.O(un1_inf_abs0_axb_13)
);
defparam \reg2_RNIKN0A[13] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIMO0A[14]  (
	.I0(inf_abs0_2[14]),
	.I1(reg2[14]),
	.O(un1_inf_abs0_axb_14)
);
defparam \reg2_RNIMO0A[14] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIOP0A[15]  (
	.I0(inf_abs0_2[15]),
	.I1(reg2[15]),
	.O(un1_inf_abs0_axb_15)
);
defparam \reg2_RNIOP0A[15] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIQQ0A[16]  (
	.I0(inf_abs0_2[16]),
	.I1(reg2[16]),
	.O(un1_inf_abs0_axb_16)
);
defparam \reg2_RNIQQ0A[16] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNISR0A[17]  (
	.I0(inf_abs0_2[17]),
	.I1(reg2[17]),
	.O(un1_inf_abs0_axb_17)
);
defparam \reg2_RNISR0A[17] .INIT=4'h6;
// @7:74
  LUT2 \reg2_RNIUS0A[18]  (
	.I0(inf_abs0_2[18]),
	.I1(reg2[18]),
	.O(un1_inf_abs0_axb_18)
);
defparam \reg2_RNIUS0A[18] .INIT=4'h6;
// @7:74
  LUT2 un1_inf_abs0_0_cry_0_RNO (
	.I0(inf_abs0_2[0]),
	.I1(reg1[0]),
	.O(un1_inf_abs0_11[0])
);
defparam un1_inf_abs0_0_cry_0_RNO.INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIDDEN[1]  (
	.I0(inf_abs0_2[1]),
	.I1(reg1[1]),
	.O(un1_inf_abs0_0_axb_1)
);
defparam \reg1_RNIDDEN[1] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIFEEN[2]  (
	.I0(inf_abs0_2[2]),
	.I1(reg1[2]),
	.O(un1_inf_abs0_0_axb_2)
);
defparam \reg1_RNIFEEN[2] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIHFEN[3]  (
	.I0(inf_abs0_2[3]),
	.I1(reg1[3]),
	.O(un1_inf_abs0_0_axb_3)
);
defparam \reg1_RNIHFEN[3] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIJGEN[4]  (
	.I0(inf_abs0_2[4]),
	.I1(reg1[4]),
	.O(un1_inf_abs0_0_axb_4)
);
defparam \reg1_RNIJGEN[4] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNILHEN[5]  (
	.I0(inf_abs0_2[5]),
	.I1(reg1[5]),
	.O(un1_inf_abs0_0_axb_5)
);
defparam \reg1_RNILHEN[5] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNINIEN[6]  (
	.I0(inf_abs0_2[6]),
	.I1(reg1[6]),
	.O(un1_inf_abs0_0_axb_6)
);
defparam \reg1_RNINIEN[6] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIPJEN[7]  (
	.I0(inf_abs0_2[7]),
	.I1(reg1[7]),
	.O(un1_inf_abs0_0_axb_7)
);
defparam \reg1_RNIPJEN[7] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIRKEN[8]  (
	.I0(inf_abs0_2[8]),
	.I1(reg1[8]),
	.O(un1_inf_abs0_0_axb_8)
);
defparam \reg1_RNIRKEN[8] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNITLEN[9]  (
	.I0(inf_abs0_2[9]),
	.I1(reg1[9]),
	.O(un1_inf_abs0_0_axb_9)
);
defparam \reg1_RNITLEN[9] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIDGQL[10]  (
	.I0(inf_abs0_2[10]),
	.I1(reg1[10]),
	.O(un1_inf_abs0_0_axb_10)
);
defparam \reg1_RNIDGQL[10] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIFHQL[11]  (
	.I0(inf_abs0_2[11]),
	.I1(reg1[11]),
	.O(un1_inf_abs0_0_axb_11)
);
defparam \reg1_RNIFHQL[11] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIHIQL[12]  (
	.I0(inf_abs0_2[12]),
	.I1(reg1[12]),
	.O(un1_inf_abs0_0_axb_12)
);
defparam \reg1_RNIHIQL[12] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIJJQL[13]  (
	.I0(inf_abs0_2[13]),
	.I1(reg1[13]),
	.O(un1_inf_abs0_0_axb_13)
);
defparam \reg1_RNIJJQL[13] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNILKQL[14]  (
	.I0(inf_abs0_2[14]),
	.I1(reg1[14]),
	.O(un1_inf_abs0_0_axb_14)
);
defparam \reg1_RNILKQL[14] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNINLQL[15]  (
	.I0(inf_abs0_2[15]),
	.I1(reg1[15]),
	.O(un1_inf_abs0_0_axb_15)
);
defparam \reg1_RNINLQL[15] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIPMQL[16]  (
	.I0(inf_abs0_2[16]),
	.I1(reg1[16]),
	.O(un1_inf_abs0_0_axb_16)
);
defparam \reg1_RNIPMQL[16] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNIRNQL[17]  (
	.I0(inf_abs0_2[17]),
	.I1(reg1[17]),
	.O(un1_inf_abs0_0_axb_17)
);
defparam \reg1_RNIRNQL[17] .INIT=4'h6;
// @7:74
  LUT2 \reg1_RNITOQL[18]  (
	.I0(inf_abs0_2[18]),
	.I1(reg1[18]),
	.O(un1_inf_abs0_0_axb_18)
);
defparam \reg1_RNITOQL[18] .INIT=4'h6;
// @7:95
  LUT1 un3_reg3_axb_1_cZ (
	.I0(reg3[4]),
	.O(un3_reg3_axb_1)
);
defparam un3_reg3_axb_1_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_2_cZ (
	.I0(reg3[5]),
	.O(un3_reg3_axb_2)
);
defparam un3_reg3_axb_2_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_3_cZ (
	.I0(reg3[6]),
	.O(un3_reg3_axb_3)
);
defparam un3_reg3_axb_3_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_4_cZ (
	.I0(reg3[7]),
	.O(un3_reg3_axb_4)
);
defparam un3_reg3_axb_4_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_5_cZ (
	.I0(reg3[8]),
	.O(un3_reg3_axb_5)
);
defparam un3_reg3_axb_5_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_6_cZ (
	.I0(reg3[9]),
	.O(un3_reg3_axb_6)
);
defparam un3_reg3_axb_6_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_7_cZ (
	.I0(reg3[10]),
	.O(un3_reg3_axb_7)
);
defparam un3_reg3_axb_7_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_8_cZ (
	.I0(reg3[11]),
	.O(un3_reg3_axb_8)
);
defparam un3_reg3_axb_8_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_9_cZ (
	.I0(reg3[12]),
	.O(un3_reg3_axb_9)
);
defparam un3_reg3_axb_9_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_10_cZ (
	.I0(reg3[13]),
	.O(un3_reg3_axb_10)
);
defparam un3_reg3_axb_10_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_11_cZ (
	.I0(reg3[14]),
	.O(un3_reg3_axb_11)
);
defparam un3_reg3_axb_11_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_12_cZ (
	.I0(reg3[15]),
	.O(un3_reg3_axb_12)
);
defparam un3_reg3_axb_12_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_13_cZ (
	.I0(reg3[16]),
	.O(un3_reg3_axb_13)
);
defparam un3_reg3_axb_13_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_14_cZ (
	.I0(reg3[17]),
	.O(un3_reg3_axb_14)
);
defparam un3_reg3_axb_14_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_15_cZ (
	.I0(reg3[18]),
	.O(un3_reg3_axb_15)
);
defparam un3_reg3_axb_15_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_16_cZ (
	.I0(reg3[19]),
	.O(un3_reg3_axb_16)
);
defparam un3_reg3_axb_16_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_17_cZ (
	.I0(reg3[20]),
	.O(un3_reg3_axb_17)
);
defparam un3_reg3_axb_17_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_18_cZ (
	.I0(reg3[21]),
	.O(un3_reg3_axb_18)
);
defparam un3_reg3_axb_18_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_19_cZ (
	.I0(reg3[22]),
	.O(un3_reg3_axb_19)
);
defparam un3_reg3_axb_19_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_20_cZ (
	.I0(reg3[23]),
	.O(un3_reg3_axb_20)
);
defparam un3_reg3_axb_20_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_21_cZ (
	.I0(reg3[24]),
	.O(un3_reg3_axb_21)
);
defparam un3_reg3_axb_21_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_22_cZ (
	.I0(reg3[25]),
	.O(un3_reg3_axb_22)
);
defparam un3_reg3_axb_22_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_23_cZ (
	.I0(reg3[26]),
	.O(un3_reg3_axb_23)
);
defparam un3_reg3_axb_23_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_24_cZ (
	.I0(reg3[27]),
	.O(un3_reg3_axb_24)
);
defparam un3_reg3_axb_24_cZ.INIT=2'h2;
// @7:95
  LUT1 un3_reg3_axb_25_cZ (
	.I0(reg3[28]),
	.O(un3_reg3_axb_25)
);
defparam un3_reg3_axb_25_cZ.INIT=2'h2;
// @7:466
  LUT1 un3_t_s_1_RNIB3TC (
	.I0(un3_t_s_1),
	.O(N_4541_i)
);
defparam un3_t_s_1_RNIB3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_2_RNIC3TC (
	.I0(un3_t_s_2),
	.O(N_4542_i)
);
defparam un3_t_s_2_RNIC3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_3_RNID3TC (
	.I0(un3_t_s_3),
	.O(N_4543_i)
);
defparam un3_t_s_3_RNID3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_4_RNIE3TC (
	.I0(un3_t_s_4),
	.O(N_4544_i)
);
defparam un3_t_s_4_RNIE3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_5_RNIF3TC (
	.I0(un3_t_s_5),
	.O(N_4545_i)
);
defparam un3_t_s_5_RNIF3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_6_RNIG3TC (
	.I0(un3_t_s_6),
	.O(N_4546_i)
);
defparam un3_t_s_6_RNIG3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_7_RNIH3TC (
	.I0(un3_t_s_7),
	.O(N_4547_i)
);
defparam un3_t_s_7_RNIH3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_8_RNII3TC (
	.I0(un3_t_s_8),
	.O(N_4548_i)
);
defparam un3_t_s_8_RNII3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_9_RNIJ3TC (
	.I0(un3_t_s_9),
	.O(N_4549_i)
);
defparam un3_t_s_9_RNIJ3TC.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_10_RNIRF0A (
	.I0(un3_t_s_10),
	.O(N_4550_i)
);
defparam un3_t_s_10_RNIRF0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_11_RNISF0A (
	.I0(un3_t_s_11),
	.O(N_4551_i)
);
defparam un3_t_s_11_RNISF0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_12_RNITF0A (
	.I0(un3_t_s_12),
	.O(N_4552_i)
);
defparam un3_t_s_12_RNITF0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_13_RNIUF0A (
	.I0(un3_t_s_13),
	.O(N_4553_i)
);
defparam un3_t_s_13_RNIUF0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_14_RNIVF0A (
	.I0(un3_t_s_14),
	.O(N_4554_i)
);
defparam un3_t_s_14_RNIVF0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_15_RNI0G0A (
	.I0(un3_t_s_15),
	.O(N_4555_i)
);
defparam un3_t_s_15_RNI0G0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_16_RNI1G0A (
	.I0(un3_t_s_16),
	.O(N_4556_i)
);
defparam un3_t_s_16_RNI1G0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_17_RNI2G0A (
	.I0(un3_t_s_17),
	.O(N_4557_i)
);
defparam un3_t_s_17_RNI2G0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_18_RNI3G0A (
	.I0(un3_t_s_18),
	.O(N_4558_i)
);
defparam un3_t_s_18_RNI3G0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_19_RNI4G0A (
	.I0(un3_t_s_19),
	.O(N_4559_i)
);
defparam un3_t_s_19_RNI4G0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_20_RNISG0A (
	.I0(un3_t_s_20),
	.O(N_4560_i)
);
defparam un3_t_s_20_RNISG0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_21_RNITG0A (
	.I0(un3_t_s_21),
	.O(N_4561_i)
);
defparam un3_t_s_21_RNITG0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_22_RNIUG0A (
	.I0(un3_t_s_22),
	.O(N_4562_i)
);
defparam un3_t_s_22_RNIUG0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_23_RNIVG0A (
	.I0(un3_t_s_23),
	.O(N_4563_i)
);
defparam un3_t_s_23_RNIVG0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_24_RNI0H0A (
	.I0(un3_t_s_24),
	.O(N_4564_i)
);
defparam un3_t_s_24_RNI0H0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_25_RNI1H0A (
	.I0(un3_t_s_25),
	.O(N_4565_i)
);
defparam un3_t_s_25_RNI1H0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_26_RNI2H0A (
	.I0(un3_t_s_26),
	.O(N_4566_i)
);
defparam un3_t_s_26_RNI2H0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_27_RNI3H0A (
	.I0(un3_t_s_27),
	.O(N_4567_i)
);
defparam un3_t_s_27_RNI3H0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_28_RNI4H0A (
	.I0(un3_t_s_28),
	.O(N_4568_i)
);
defparam un3_t_s_28_RNI4H0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_29_RNI5H0A (
	.I0(un3_t_s_29),
	.O(N_4569_i)
);
defparam un3_t_s_29_RNI5H0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_30_RNITH0A (
	.I0(un3_t_s_30),
	.O(N_4570_i)
);
defparam un3_t_s_30_RNITH0A.INIT=2'h1;
// @7:466
  LUT1 un3_t_s_31_RNIUH0A (
	.I0(un3_t_s_31),
	.O(N_4571_i)
);
defparam un3_t_s_31_RNIUH0A.INIT=2'h1;
// @7:83
  LUT2 inf_abs0_2_axb_29_cZ (
	.I0(ir[29]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_29)
);
defparam inf_abs0_2_axb_29_cZ.INIT=4'h6;
// @7:151
  LUT4 un26_r_df30_cZ (
	.I0(m_2[30]),
	.I1(m_2_i[31]),
	.I2(r_4_i[31]),
	.I3(r_6[30]),
	.O(un26_r_df30)
);
defparam un26_r_df30_cZ.INIT=16'h8241;
// @7:128
  LUT4 \d_cnst_sn.un14_r_0_I_88  (
	.I0(m_2[30]),
	.I1(m_2[31]),
	.I2(r_4[30]),
	.I3(r_4[31]),
	.O(un14_r_0_N_2)
);
defparam \d_cnst_sn.un14_r_0_I_88 .INIT=16'h8421;
// @7:47
  FDC b_Z (
	.Q(b),
	.D(b_0),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDCE \d_Z[0]  (
	.Q(d[0]),
	.D(d_cnst[0]),
	.C(clock),
	.CLR(reset),
	.CE(dce[0])
);
// @7:47
  FDCE \d_Z[1]  (
	.Q(d[1]),
	.D(d_cnst_sm0),
	.C(clock),
	.CLR(reset),
	.CE(dce[0])
);
// @7:47
  FDC \ir_Z[22]  (
	.Q(ir[22]),
	.D(ir_3[22]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[23]  (
	.Q(ir[23]),
	.D(ir_3[23]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[24]  (
	.Q(ir[24]),
	.D(ir_3[24]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[25]  (
	.Q(ir[25]),
	.D(ir_3[25]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[26]  (
	.Q(ir[26]),
	.D(ir_3[26]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[27]  (
	.Q(ir[27]),
	.D(ir_3[27]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[28]  (
	.Q(ir[28]),
	.D(ir_3[28]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[29]  (
	.Q(ir[29]),
	.D(ir_3[29]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[30]  (
	.Q(ir[30]),
	.D(ir_3[30]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[31]  (
	.Q(ir[31]),
	.D(ir_3[31]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[7]  (
	.Q(ir[7]),
	.D(ir_3[7]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[8]  (
	.Q(ir[8]),
	.D(ir_3[8]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[9]  (
	.Q(ir[9]),
	.D(ir_3[9]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[10]  (
	.Q(ir[10]),
	.D(ir_3[10]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[11]  (
	.Q(ir[11]),
	.D(ir_3[11]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[12]  (
	.Q(ir[12]),
	.D(ir_3[12]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[13]  (
	.Q(ir[13]),
	.D(ir_3[13]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[14]  (
	.Q(ir[14]),
	.D(ir_3[14]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[15]  (
	.Q(ir[15]),
	.D(ir_3[15]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[16]  (
	.Q(ir[16]),
	.D(ir_3[16]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[17]  (
	.Q(ir[17]),
	.D(ir_3[17]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[18]  (
	.Q(ir[18]),
	.D(ir_3[18]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[19]  (
	.Q(ir[19]),
	.D(ir_3[19]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[20]  (
	.Q(ir[20]),
	.D(ir_3[20]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[21]  (
	.Q(ir[21]),
	.D(ir_3[21]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[0]  (
	.Q(ir[0]),
	.D(ir_3[0]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[1]  (
	.Q(ir[1]),
	.D(ir_3[1]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[2]  (
	.Q(ir[2]),
	.D(ir_3[2]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[3]  (
	.Q(ir[3]),
	.D(ir_3[3]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[4]  (
	.Q(ir[4]),
	.D(ir_3[4]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[5]  (
	.Q(ir[5]),
	.D(ir_3[5]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_Z[6]  (
	.Q(ir[6]),
	.D(ir_3[6]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDCE \reg0_Z[31]  (
	.Q(reg0[31]),
	.D(N_3856_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[16]  (
	.Q(reg0[16]),
	.D(reg0_28[16]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[17]  (
	.Q(reg0[17]),
	.D(reg0_28[17]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[18]  (
	.Q(reg0[18]),
	.D(reg0_28[18]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[19]  (
	.Q(reg0[19]),
	.D(N_3829_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[20]  (
	.Q(reg0[20]),
	.D(N_3803_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[21]  (
	.Q(reg0[21]),
	.D(N_3777_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[22]  (
	.Q(reg0[22]),
	.D(N_3751_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[23]  (
	.Q(reg0[23]),
	.D(N_3725_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[24]  (
	.Q(reg0[24]),
	.D(N_3699_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[25]  (
	.Q(reg0[25]),
	.D(N_3673_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[26]  (
	.Q(reg0[26]),
	.D(N_3341_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[27]  (
	.Q(reg0[27]),
	.D(N_3315_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[28]  (
	.Q(reg0[28]),
	.D(N_3289_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[29]  (
	.Q(reg0[29]),
	.D(N_3569_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[30]  (
	.Q(reg0[30]),
	.D(N_3550_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[1]  (
	.Q(reg0[1]),
	.D(reg0_28[1]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[2]  (
	.Q(reg0[2]),
	.D(reg0_28[2]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[3]  (
	.Q(reg0[3]),
	.D(reg0_28[3]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[4]  (
	.Q(reg0[4]),
	.D(reg0_28[4]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[5]  (
	.Q(reg0[5]),
	.D(reg0_28[5]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[6]  (
	.Q(reg0[6]),
	.D(reg0_28[6]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[7]  (
	.Q(reg0[7]),
	.D(reg0_28_7_rep1),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[8]  (
	.Q(reg0[8]),
	.D(reg0_28[8]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[9]  (
	.Q(reg0[9]),
	.D(reg0_28[9]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[10]  (
	.Q(reg0[10]),
	.D(reg0_28[10]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[11]  (
	.Q(reg0[11]),
	.D(reg0_28[11]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[12]  (
	.Q(reg0[12]),
	.D(reg0_28[12]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[13]  (
	.Q(reg0[13]),
	.D(reg0_28[13]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[14]  (
	.Q(reg0[14]),
	.D(reg0_28[14]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg0_Z[15]  (
	.Q(reg0[15]),
	.D(reg0_28[15]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg1_Z[18]  (
	.Q(reg1[18]),
	.D(reg1_16[18]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[19]  (
	.Q(reg1[19]),
	.D(reg0_28_3_2492),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[20]  (
	.Q(reg1[20]),
	.D(reg0_28_4_2459),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[21]  (
	.Q(reg1[21]),
	.D(reg0_28_5_2426),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[22]  (
	.Q(reg1[22]),
	.D(reg0_28_6_2393),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[23]  (
	.Q(reg1[23]),
	.D(reg0_28_7_2360),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[24]  (
	.Q(reg1[24]),
	.D(reg0_28_8_2327),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[25]  (
	.Q(reg1[25]),
	.D(N_3673),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[26]  (
	.Q(reg1[26]),
	.D(reg1_16_7_1870),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[27]  (
	.Q(reg1[27]),
	.D(reg1_16_8_1837),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[28]  (
	.Q(reg1[28]),
	.D(reg1_16_9),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[29]  (
	.Q(reg1[29]),
	.D(reg0_28_10_2261_a6_3_2_lut6_2_RNIOK9O5),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[30]  (
	.Q(reg1[30]),
	.D(N_3550),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[31]  (
	.Q(reg1[31]),
	.D(N_3856),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg0_Z[0]  (
	.Q(reg0[0]),
	.D(reg0_28[0]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_4_i)
);
// @7:47
  FDCE \reg1_Z[3]  (
	.Q(reg1[3]),
	.D(reg1_16[3]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[4]  (
	.Q(reg1[4]),
	.D(reg1_16[4]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[5]  (
	.Q(reg1[5]),
	.D(reg1_16[5]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[6]  (
	.Q(reg1[6]),
	.D(reg1_16[6]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[7]  (
	.Q(reg1[7]),
	.D(reg0_28[7]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[8]  (
	.Q(reg1[8]),
	.D(reg1_16[8]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[9]  (
	.Q(reg1[9]),
	.D(reg1_16[9]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[10]  (
	.Q(reg1[10]),
	.D(reg1_16[10]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[11]  (
	.Q(reg1[11]),
	.D(reg1_16[11]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[12]  (
	.Q(reg1[12]),
	.D(reg1_16[12]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[13]  (
	.Q(reg1[13]),
	.D(reg1_16[13]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[14]  (
	.Q(reg1[14]),
	.D(reg1_16[14]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[15]  (
	.Q(reg1[15]),
	.D(reg1_16[15]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[16]  (
	.Q(reg1[16]),
	.D(reg1_16[16]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[17]  (
	.Q(reg1[17]),
	.D(reg1_16[17]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg2_Z[20]  (
	.Q(reg2[20]),
	.D(reg2_16[20]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[21]  (
	.Q(reg2[21]),
	.D(reg2_16[21]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[22]  (
	.Q(reg2[22]),
	.D(reg2_16[22]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[23]  (
	.Q(reg2[23]),
	.D(reg2_16[23]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[24]  (
	.Q(reg2[24]),
	.D(reg2_16[24]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[25]  (
	.Q(reg2[25]),
	.D(reg2_16[25]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[26]  (
	.Q(reg2[26]),
	.D(reg2_16[26]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[27]  (
	.Q(reg2[27]),
	.D(reg2_16[27]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[28]  (
	.Q(reg2[28]),
	.D(reg2_16[28]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[29]  (
	.Q(reg2[29]),
	.D(reg2_16[29]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[30]  (
	.Q(reg2[30]),
	.D(reg2_16[30]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[31]  (
	.Q(reg2[31]),
	.D(reg2_16[31]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg1_Z[0]  (
	.Q(reg1[0]),
	.D(reg1_16[0]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[1]  (
	.Q(reg1[1]),
	.D(reg1_16[1]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg1_Z[2]  (
	.Q(reg1[2]),
	.D(reg1_16[2]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_3_i)
);
// @7:47
  FDCE \reg2_Z[5]  (
	.Q(reg2[5]),
	.D(reg2_16[5]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[6]  (
	.Q(reg2[6]),
	.D(reg2_16[6]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[7]  (
	.Q(reg2[7]),
	.D(reg2_16[7]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[8]  (
	.Q(reg2[8]),
	.D(reg2_16[8]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[9]  (
	.Q(reg2[9]),
	.D(reg2_16[9]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[10]  (
	.Q(reg2[10]),
	.D(reg2_16[10]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[11]  (
	.Q(reg2[11]),
	.D(reg2_16[11]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[12]  (
	.Q(reg2[12]),
	.D(reg2_16[12]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[13]  (
	.Q(reg2[13]),
	.D(reg2_16[13]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[14]  (
	.Q(reg2[14]),
	.D(reg2_16[14]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[15]  (
	.Q(reg2[15]),
	.D(reg2_16[15]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[16]  (
	.Q(reg2[16]),
	.D(reg2_16[16]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[17]  (
	.Q(reg2[17]),
	.D(reg2_16[17]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[18]  (
	.Q(reg2[18]),
	.D(reg2_16[18]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[19]  (
	.Q(reg2[19]),
	.D(reg2_16[19]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \datao_Z[22]  (
	.Q(datao[22]),
	.D(r_4_3_1690_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[23]  (
	.Q(datao[23]),
	.D(r_4_3_0_1664_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[24]  (
	.Q(datao[24]),
	.D(r_4_3_1_1638_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[25]  (
	.Q(datao[25]),
	.D(r_4_3_2_1612_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[26]  (
	.Q(datao[26]),
	.D(r_4_3_3_1586_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[27]  (
	.Q(datao[27]),
	.D(r_4_3_4_1560_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[28]  (
	.Q(datao[28]),
	.D(r_4_3_5_1534_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[29]  (
	.Q(datao[29]),
	.D(r_4_3_6_1508_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[30]  (
	.Q(datao[30]),
	.D(r_4_3_lut6_2_O5[30]),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[31]  (
	.Q(datao[31]),
	.D(r_4_3_8_1467),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \reg2_Z[0]  (
	.Q(reg2[0]),
	.D(reg2_16[0]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[1]  (
	.Q(reg2[1]),
	.D(reg2_16[1]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[2]  (
	.Q(reg2[2]),
	.D(reg2_16[2]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[3]  (
	.Q(reg2[3]),
	.D(reg2_16[3]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \reg2_Z[4]  (
	.Q(reg2[4]),
	.D(reg2_16[4]),
	.C(clock),
	.CLR(reset),
	.CE(un1_state_1_0_i)
);
// @7:47
  FDCE \datao_Z[7]  (
	.Q(datao[7]),
	.D(r_4_3_9_1442_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[8]  (
	.Q(datao[8]),
	.D(r_4_3_10_1416_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[9]  (
	.Q(datao[9]),
	.D(r_4_3_11_1390_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[10]  (
	.Q(datao[10]),
	.D(r_4_3_12_1364_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[11]  (
	.Q(datao[11]),
	.D(r_4_3_13_1338_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[12]  (
	.Q(datao[12]),
	.D(r_4_3_14_1312_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[13]  (
	.Q(datao[13]),
	.D(r_4_3_15_1286_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[14]  (
	.Q(datao[14]),
	.D(r_4_3_16_1260_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[15]  (
	.Q(datao[15]),
	.D(r_4_3_17_1234_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[16]  (
	.Q(datao[16]),
	.D(r_4_3_18_1208_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[17]  (
	.Q(datao[17]),
	.D(r_4_3_19_1182_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[18]  (
	.Q(datao[18]),
	.D(r_4_3_20_1156_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[19]  (
	.Q(datao[19]),
	.D(N_2724),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[20]  (
	.Q(datao[20]),
	.D(r_4_3_22_1104_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[21]  (
	.Q(datao[21]),
	.D(r_4_3_23_1078_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \addr_Z[12]  (
	.Q(addr[12]),
	.D(N_2656_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[13]  (
	.Q(addr[13]),
	.D(N_2636_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[14]  (
	.Q(addr[14]),
	.D(N_2616_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[15]  (
	.Q(addr[15]),
	.D(N_2596_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[16]  (
	.Q(addr[16]),
	.D(N_2576_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[17]  (
	.Q(addr[17]),
	.D(N_2556_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[18]  (
	.Q(addr[18]),
	.D(N_2536_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[19]  (
	.Q(addr[19]),
	.D(N_2516_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \datao_Z[0]  (
	.Q(datao[0]),
	.D(r_4_3_24_836_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[1]  (
	.Q(datao[1]),
	.D(r_4_3_25_810_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[2]  (
	.Q(datao[2]),
	.D(N_36_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[3]  (
	.Q(datao[3]),
	.D(r_4_3_27_758_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[4]  (
	.Q(datao[4]),
	.D(r_4_3_28_732_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[5]  (
	.Q(datao[5]),
	.D(r_4_3_29_706_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \datao_Z[6]  (
	.Q(datao[6]),
	.D(r_4_3_30_680_i_m2),
	.C(clock),
	.CLR(reset),
	.CE(addr_4_sqmuxa_1)
);
// @7:47
  FDCE \reg3_Z[26]  (
	.Q(reg3[26]),
	.D(reg3_17[26]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[27]  (
	.Q(reg3[27]),
	.D(reg3_17[27]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[28]  (
	.Q(reg3[28]),
	.D(reg3_17[28]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \addr_Z[0]  (
	.Q(addr[0]),
	.D(N_2335_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[1]  (
	.Q(addr[1]),
	.D(N_2315_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[2]  (
	.Q(addr[2]),
	.D(N_47_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[3]  (
	.Q(addr[3]),
	.D(N_2267_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[4]  (
	.Q(addr[4]),
	.D(N_56_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[5]  (
	.Q(addr[5]),
	.D(N_2219_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[6]  (
	.Q(addr[6]),
	.D(N_2199_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[7]  (
	.Q(addr[7]),
	.D(N_2179_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[8]  (
	.Q(addr[8]),
	.D(N_2159_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[9]  (
	.Q(addr[9]),
	.D(N_2139_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[10]  (
	.Q(addr[10]),
	.D(N_2119_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \addr_Z[11]  (
	.Q(addr[11]),
	.D(N_2099_i),
	.C(clock),
	.CLR(reset),
	.CE(addr_0_sqmuxa_1_i)
);
// @7:47
  FDCE \reg3_Z[11]  (
	.Q(reg3[11]),
	.D(reg3_17[11]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[12]  (
	.Q(reg3[12]),
	.D(reg3_17[12]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[13]  (
	.Q(reg3[13]),
	.D(reg3_17[13]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[14]  (
	.Q(reg3[14]),
	.D(reg3_17[14]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[15]  (
	.Q(reg3[15]),
	.D(reg3_17[15]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[16]  (
	.Q(reg3[16]),
	.D(reg3_17[16]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[17]  (
	.Q(reg3[17]),
	.D(reg3_17[17]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[18]  (
	.Q(reg3[18]),
	.D(reg3_17[18]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[19]  (
	.Q(reg3[19]),
	.D(reg3_17[19]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[20]  (
	.Q(reg3[20]),
	.D(reg3_17[20]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[21]  (
	.Q(reg3[21]),
	.D(reg3_17[21]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[22]  (
	.Q(reg3[22]),
	.D(reg3_17[22]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[23]  (
	.Q(reg3[23]),
	.D(reg3_17[23]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[24]  (
	.Q(reg3[24]),
	.D(reg3_17[24]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[25]  (
	.Q(reg3[25]),
	.D(reg3_17[25]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[0]  (
	.Q(reg3[0]),
	.D(reg3_17[0]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[1]  (
	.Q(reg3[1]),
	.D(reg3_17[1]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[2]  (
	.Q(reg3[2]),
	.D(reg3_17[2]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[3]  (
	.Q(reg3[3]),
	.D(\d_cnst_sn.reg3_N_7_i ),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[4]  (
	.Q(reg3[4]),
	.D(reg3_17[4]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[5]  (
	.Q(reg3[5]),
	.D(reg3_17[5]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[6]  (
	.Q(reg3[6]),
	.D(reg3_17[6]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[7]  (
	.Q(reg3[7]),
	.D(reg3_17[7]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[8]  (
	.Q(reg3[8]),
	.D(reg3_17[8]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[9]  (
	.Q(reg3[9]),
	.D(reg3_17[9]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDCE \reg3_Z[10]  (
	.Q(reg3[10]),
	.D(reg3_17[10]),
	.C(clock),
	.CLR(reset),
	.CE(state[0])
);
// @7:47
  FDC rd_Z (
	.Q(rd),
	.D(rd_18),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \state_Z[0]  (
	.Q(state[0]),
	.D(state_i[0]),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC wr_Z (
	.Q(wr),
	.D(addr_4_sqmuxa_1),
	.C(clock),
	.CLR(reset)
);
// @7:47
  FDC \ir_fast_Z[31]  (
	.Q(ir_fast[31]),
	.D(ir_3_fast[31]),
	.C(clock),
	.CLR(reset)
);
// @7:83
  MUXCY_L inf_abs0_2_cry_29_outext (
	.DI(GND),
	.CI(inf_abs0_2_cry_29_0),
	.S(inf_abs0_2_cry_29_1),
	.LO(inf_abs0_2_cry_29)
);
// @7:95
  MUXCY un3_reg3_cry_25_outext (
	.DI(GND),
	.CI(un3_reg3_cry_25_0),
	.S(un3_reg3_cry_25_1),
	.O(un3_reg3_cry_25)
);
// @7:83
  MUXCY inf_abs0_2_cry_30_outext (
	.DI(GND),
	.CI(inf_abs0_2_0[31]),
	.S(inf_abs0_2_1[31]),
	.O(inf_abs0_2[31])
);
// @7:128
  MUXCY un14_r_0_I_83_cZ (
	.DI(GND),
	.CI(un14_r_0_data_tmp[9]),
	.S(un14_r_0_N_2),
	.O(un14_r_0_I_83)
);
// @7:118
  MUXCY \un11_r_cry_cZ[30]  (
	.DI(un11_r_lt30),
	.CI(un11_r_cry[28]),
	.S(un11_r_df30),
	.O(un11_r_cry[30])
);
// @7:143
  MUXCY \b18_cry[30]  (
	.DI(b18_lt30),
	.CI(b18_cry[28]),
	.S(b18_df30),
	.O(b18)
);
// @7:151
  MUXCY \un26_r_cry_cZ[30]  (
	.DI(un26_r_lt30),
	.CI(un26_r_cry[28]),
	.S(un26_r_df30),
	.O(un26_r_cry[30])
);
// @7:83
  MUXCY inf_abs0_2_cry_29_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_28),
	.S(inf_abs0_2_axb_29),
	.O(inf_abs0_2_cry_29_0)
);
// @7:246
  LUT5 \d_cnst_sn.un87_df  (
	.I0(d[0]),
	.I1(d[1]),
	.I2(d_cnst_ss0_x),
	.I3(un1_df_1),
	.I4(d_cnst_sm0),
	.O(un87_df)
);
defparam \d_cnst_sn.un87_df .INIT=32'h88F08800;
// @7:47
  LUT4_L \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_RNIOK9O5  (
	.I0(\d_cnst_sn.g0_0_2 ),
	.I1(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I2(t_1[29]),
	.I3(\d_cnst_sn.g0_rn_1 ),
	.LO(reg0_28_10_2261_a6_3_2_lut6_2_RNIOK9O5)
);
defparam \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_RNIOK9O5 .INIT=16'hFF02;
// @7:103
  LUT6 \d_cnst_sn.un1_cf_x_RNI07TU1  (
	.I0(inf_abs0_2[23]),
	.I1(un36_df),
	.I2(N_1890),
	.I3(m7),
	.I4(un1_cf_x),
	.I5(un87_df),
	.O(\d_cnst_sn.reg3_17_sn_m7_0 )
);
defparam \d_cnst_sn.un1_cf_x_RNI07TU1 .INIT=64'h0000FFFEFFFEFFFE;
// @7:103
  LUT4 \d_cnst_sn.un1_cf_x  (
	.I0(inf_abs0_2[23]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(\d_cnst_sn.reg3_5_sqmuxa_2_1 ),
	.O(un1_cf_x)
);
defparam \d_cnst_sn.un1_cf_x .INIT=16'h0400;
// @7:213
  LUT3 \d_cnst_sn.d_cnst_ss0_x  (
	.I0(inf_abs0_2[24]),
	.I1(inf_abs0_2[25]),
	.I2(inf_abs0_2[26]),
	.O(d_cnst_ss0_x)
);
defparam \d_cnst_sn.d_cnst_ss0_x .INIT=8'hBA;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNI0TVT3[7]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg0_1 [7]),
	.I4(t_1[7]),
	.I5(N_1042),
	.LO(reg0_28_7_rep1)
);
defparam \d_cnst_sn.reg0_28_6_RNI0TVT3[7] .INIT=64'h0F00FF0001001100;
// @7:358
  LUT6 \d_cnst_sn.m_2_i[0]  (
	.I0(datai[0]),
	.I1(inf_abs0_2_axb_30),
	.I2(inf_abs0_2[0]),
	.I3(inf_abs0_2_cry_29),
	.I4(inf_abs0_2[27]),
	.I5(inf_abs0_2[28]),
	.O(m_2_i[0])
);
defparam \d_cnst_sn.m_2_i[0] .INIT=64'h1D551D551D550F0F;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_RNIC3O74  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.g0_1 ),
	.I3(un32_reg0_s_29),
	.I4(un11_reg0_s_29),
	.LO(\d_cnst_sn.g0_rn_1 )
);
defparam \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_RNIC3O74 .INIT=32'hFAF8F2F0;
// @7:213
  LUT6 \d_cnst_sn.un1_df_1  (
	.I0(b),
	.I1(inf_abs0_2_axb_30),
	.I2(inf_abs0_2_cry_29),
	.I3(inf_abs0_2[24]),
	.I4(inf_abs0_2[25]),
	.I5(inf_abs0_2[26]),
	.O(un1_df_1)
);
defparam \d_cnst_sn.un1_df_1 .INIT=64'h2A3F2A1500000000;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_RNIQARE5  (
	.I0(\d_cnst_sn.g0_0_2 ),
	.I1(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I2(\d_cnst_sn.g0_1 ),
	.I3(t_1[29]),
	.I4(\d_cnst_sn.g3 ),
	.LO(N_3569_rep1)
);
defparam \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_RNIQARE5 .INIT=32'hFCFEF0F2;
// @7:47
  LUT6_L \d_cnst_sn.reg0_28_3_2492_rep1  (
	.I0(\d_cnst_sn.reg0_28_2526_a5_1_0 ),
	.I1(\d_cnst_sn.reg1_16_8_1837_2_tz ),
	.I2(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I3(\d_cnst_sn.reg0_28_0 [19]),
	.I4(t_1[19]),
	.I5(\d_cnst_sn.reg0_28_3_2492_1 ),
	.LO(N_3829_rep1)
);
defparam \d_cnst_sn.reg0_28_3_2492_rep1 .INIT=64'hFFFFFFFF0E00EE00;
// @7:47
  LUT6_L \d_cnst_sn.reg0_28_4_2459_rep1  (
	.I0(\d_cnst_sn.reg0_28_2526_a5_1_0 ),
	.I1(\d_cnst_sn.reg1_16_8_1837_2_tz ),
	.I2(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I3(\d_cnst_sn.reg0_28_0 [20]),
	.I4(t_1[20]),
	.I5(\d_cnst_sn.reg0_28_4_2459_0 ),
	.LO(N_3803_rep1)
);
defparam \d_cnst_sn.reg0_28_4_2459_rep1 .INIT=64'hFFFFFFFF0E00EE00;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_5_2426_rep1  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_5_2426_3_1 ),
	.I2(\d_cnst_sn.reg0_28_5_2426_a6_1_1 ),
	.I3(t_1[21]),
	.I4(\d_cnst_sn.reg0_28_5_2426_0 ),
	.LO(N_3777_rep1)
);
defparam \d_cnst_sn.reg0_28_5_2426_rep1 .INIT=32'hFFFF54FC;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_6_2393_rep1  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_6_2393_3_1 ),
	.I2(\d_cnst_sn.reg0_28_6_2393_a6_1_1 ),
	.I3(t_1[22]),
	.I4(\d_cnst_sn.reg0_28_6_2393_0 ),
	.LO(N_3751_rep1)
);
defparam \d_cnst_sn.reg0_28_6_2393_rep1 .INIT=32'hFFFF54FC;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_7_2360_rep1  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_7_2360_3_1 ),
	.I2(\d_cnst_sn.reg0_28_7_2360_a6_1_1 ),
	.I3(t_1[23]),
	.I4(\d_cnst_sn.reg0_28_7_2360_0 ),
	.LO(N_3725_rep1)
);
defparam \d_cnst_sn.reg0_28_7_2360_rep1 .INIT=32'hFFFF54FC;
// @7:47
  LUT6_L \d_cnst_sn.reg0_28_8_2327_rep1  (
	.I0(\d_cnst_sn.reg1_16_8_1837_2_tz ),
	.I1(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I2(reg0_28_7_d[24]),
	.I3(\d_cnst_sn.reg0_28_8_2327_a6_1_1 ),
	.I4(t_1[24]),
	.I5(\d_cnst_sn.reg0_28_8_2327_0 ),
	.LO(N_3699_rep1)
);
defparam \d_cnst_sn.reg0_28_8_2327_rep1 .INIT=64'hFFFFFFFF3320FFA8;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_9_2294_rep1  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_9_2294_3_1 ),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_1_1 ),
	.I3(t_1[25]),
	.I4(\d_cnst_sn.reg0_28_9_2294_0 ),
	.LO(N_3673_rep1)
);
defparam \d_cnst_sn.reg0_28_9_2294_rep1 .INIT=32'hFFFF54FC;
// @7:47
  LUT5_L \d_cnst_sn.reg1_16_7_1870_rep1  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_10_2261_a6_1_1 ),
	.I2(\d_cnst_sn.reg1_16_7_1870_3_1 ),
	.I3(t_1[26]),
	.I4(\d_cnst_sn.reg1_16_7_1870_0 ),
	.LO(N_3341_rep1)
);
defparam \d_cnst_sn.reg1_16_7_1870_rep1 .INIT=32'hFFFF54FC;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_14_rep1  (
	.I0(inf_abs0_2[31]),
	.I1(\d_cnst_sn.reg0_28_14_2135_1_a0_2 ),
	.I2(reg3_1_1[30]),
	.I3(\d_cnst_sn.reg0_28_14_0 ),
	.I4(t_1[30]),
	.LO(N_3550_rep1)
);
defparam \d_cnst_sn.reg0_28_14_rep1 .INIT=32'hFFA0FFEC;
// @7:47
  LUT5_L \d_cnst_sn.reg1_16_8_1837_rep1  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_11_2228_a6_1_1 ),
	.I2(\d_cnst_sn.reg1_16_8_1837_3_1 ),
	.I3(t_1[27]),
	.I4(\d_cnst_sn.reg1_16_8_1837_0 ),
	.LO(N_3315_rep1)
);
defparam \d_cnst_sn.reg1_16_8_1837_rep1 .INIT=32'hFFFF54FC;
// @7:47
  LUT6_L \d_cnst_sn.reg1_16_9_rep1  (
	.I0(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I1(m_2[28]),
	.I2(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I3(\d_cnst_sn.reg1_16_9_1804_3_tz ),
	.I4(t_1[28]),
	.I5(N_3614),
	.LO(N_3289_rep1)
);
defparam \d_cnst_sn.reg1_16_9_rep1 .INIT=64'hFFFFFFFF8F88FF88;
// @7:47
  LUT6_L \d_cnst_sn.reg0_28_a1_1_lut6_2_RNIDLFQ4_0[7]  (
	.I0(b),
	.I1(inf_abs0_2[27]),
	.I2(\d_cnst_sn.g0_3_a2_2 ),
	.I3(\d_cnst_sn.g0_3_1 ),
	.I4(t_1[31]),
	.I5(t_1[30]),
	.LO(N_3856_rep1)
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_RNIDLFQ4_0[7] .INIT=64'hFF00FF30FF40FF70;
// @7:74
  LUT6 \d_cnst_sn.g0_0_0_a5_0  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(\d_cnst_sn.g0_0_0_a5_0_0 ),
	.O(N_7_0)
);
defparam \d_cnst_sn.g0_0_0_a5_0 .INIT=64'h0101010000000000;
  LUT6 \d_cnst_sn.reg0_28_a2_0_lut6_2_RNI9RAM3[2]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[31]),
	.I3(N_7_0),
	.I4(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I5(reg3_1_1[31]),
	.O(\d_cnst_sn.g0_0_0_1 )
);
defparam \d_cnst_sn.reg0_28_a2_0_lut6_2_RNI9RAM3[2] .INIT=64'hFFF1FF00FF00FF00;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_10_2261_a6_1_0_lut6_2_RNI3B3R4  (
	.I0(b),
	.I1(inf_abs0_2[27]),
	.I2(\d_cnst_sn.g0_0_0_a5_2 ),
	.I3(\d_cnst_sn.g0_0_0_1 ),
	.I4(t_1[31]),
	.I5(t_1[30]),
	.LO(reg2_16[31])
);
defparam \d_cnst_sn.reg0_28_10_2261_a6_1_0_lut6_2_RNI3B3R4 .INIT=64'hFF00FF30FF40FF70;
// @7:47
  LUT3_L \d_cnst_sn.g3_cZ  (
	.I0(N_1033),
	.I1(un32_reg0_s_29),
	.I2(un11_reg0_s_29),
	.LO(\d_cnst_sn.g3 )
);
defparam \d_cnst_sn.g3_cZ .INIT=8'hE4;
  LUT5 \d_cnst_sn.g0_0_2_cZ  (
	.I0(b),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(\d_cnst_sn.g0_0_2 )
);
defparam \d_cnst_sn.g0_0_2_cZ .INIT=32'h0000040C;
  LUT6 \d_cnst_sn.reg0_m9_i_a1_RNI2ROG2  (
	.I0(\d_cnst_sn.reg0_N_13_0 ),
	.I1(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I2(N_513_i),
	.I3(m_2[29]),
	.I4(reg0_m9_i_a1),
	.I5(reg3_1_1[29]),
	.O(\d_cnst_sn.g0_1 )
);
defparam \d_cnst_sn.reg0_m9_i_a1_RNI2ROG2 .INIT=64'hFFFFCD05FFFFCC00;
// @7:47
  LUT6 \d_cnst_sn.g0_3_a2_0  (
	.I0(datai[31]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.I5(N_7),
	.O(N_12)
);
defparam \d_cnst_sn.g0_3_a2_0 .INIT=64'h0000000800000000;
  LUT6 \d_cnst_sn.g0_3_1_cZ  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(N_12),
	.I5(reg3_1_1[31]),
	.O(\d_cnst_sn.g0_3_1 )
);
defparam \d_cnst_sn.g0_3_1_cZ .INIT=64'hFFFFFF01FFFF0000;
// @7:47
  LUT6_L \d_cnst_sn.reg0_28_a1_1_lut6_2_RNIDLFQ4[7]  (
	.I0(b),
	.I1(inf_abs0_2[27]),
	.I2(\d_cnst_sn.g0_3_a2_2 ),
	.I3(\d_cnst_sn.g0_3_1 ),
	.I4(t_1[31]),
	.I5(t_1[30]),
	.LO(N_3856)
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_RNIDLFQ4[7] .INIT=64'hFF00FF30FF40FF70;
// @7:103
  LUT4 \d_cnst_sn.reg3_17_0[28]  (
	.I0(datai[28]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_cf),
	.O(N_1685)
);
defparam \d_cnst_sn.reg3_17_0[28] .INIT=16'hA8AA;
// @7:103
  LUT4 \d_cnst_sn.reg3_17_0[27]  (
	.I0(datai[27]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_cf),
	.O(N_1684)
);
defparam \d_cnst_sn.reg3_17_0[27] .INIT=16'hA8AA;
// @7:103
  LUT4 \d_cnst_sn.reg3_17_0[26]  (
	.I0(datai[26]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_cf),
	.O(N_1683)
);
defparam \d_cnst_sn.reg3_17_0[26] .INIT=16'hA8AA;
// @7:103
  LUT4 \d_cnst_sn.reg3_17_0[25]  (
	.I0(datai[25]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_cf),
	.O(N_1682)
);
defparam \d_cnst_sn.reg3_17_0[25] .INIT=16'hA8AA;
// @7:103
  LUT4_L \d_cnst_sn.reg3_17_0[24]  (
	.I0(datai[24]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_cf),
	.LO(N_1681)
);
defparam \d_cnst_sn.reg3_17_0[24] .INIT=16'hA8AA;
// @7:103
  LUT4_L \d_cnst_sn.reg3_17_0[23]  (
	.I0(datai[23]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_cf),
	.LO(N_1680)
);
defparam \d_cnst_sn.reg3_17_0[23] .INIT=16'hA8AA;
// @7:103
  LUT4_L \d_cnst_sn.reg3_17_0[22]  (
	.I0(datai[22]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_cf),
	.LO(N_1679)
);
defparam \d_cnst_sn.reg3_17_0[22] .INIT=16'hA8AA;
// @7:103
  LUT4 \d_cnst_sn.reg3_17_0[20]  (
	.I0(datai[20]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_cf),
	.O(N_1677)
);
defparam \d_cnst_sn.reg3_17_0[20] .INIT=16'hA8AA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[7]  (
	.I0(datai[7]),
	.I1(inf_abs0_2[7]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1664)
);
defparam \d_cnst_sn.reg3_17_0[7] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[6]  (
	.I0(datai[6]),
	.I1(inf_abs0_2[6]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1663)
);
defparam \d_cnst_sn.reg3_17_0[6] .INIT=32'hAAACAAAA;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_0[2]  (
	.I0(datai[2]),
	.I1(inf_abs0_2[2]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.LO(N_1659)
);
defparam \d_cnst_sn.reg3_17_0[2] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[9]  (
	.I0(datai[9]),
	.I1(inf_abs0_2[9]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1666)
);
defparam \d_cnst_sn.reg3_17_0[9] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[11]  (
	.I0(datai[11]),
	.I1(inf_abs0_2[11]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1668)
);
defparam \d_cnst_sn.reg3_17_0[11] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[10]  (
	.I0(datai[10]),
	.I1(inf_abs0_2[10]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1667)
);
defparam \d_cnst_sn.reg3_17_0[10] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[17]  (
	.I0(datai[17]),
	.I1(inf_abs0_2[17]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1674)
);
defparam \d_cnst_sn.reg3_17_0[17] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[12]  (
	.I0(datai[12]),
	.I1(inf_abs0_2[12]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1669)
);
defparam \d_cnst_sn.reg3_17_0[12] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[18]  (
	.I0(datai[18]),
	.I1(inf_abs0_2[18]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1675)
);
defparam \d_cnst_sn.reg3_17_0[18] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[14]  (
	.I0(datai[14]),
	.I1(inf_abs0_2[14]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1671)
);
defparam \d_cnst_sn.reg3_17_0[14] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[19]  (
	.I0(datai[19]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1676)
);
defparam \d_cnst_sn.reg3_17_0[19] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[13]  (
	.I0(datai[13]),
	.I1(inf_abs0_2[13]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1670)
);
defparam \d_cnst_sn.reg3_17_0[13] .INIT=32'hAAACAAAA;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_0[1]  (
	.I0(datai[1]),
	.I1(inf_abs0_2[1]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.LO(N_1658)
);
defparam \d_cnst_sn.reg3_17_0[1] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[16]  (
	.I0(datai[16]),
	.I1(inf_abs0_2[16]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1673)
);
defparam \d_cnst_sn.reg3_17_0[16] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[15]  (
	.I0(datai[15]),
	.I1(inf_abs0_2[15]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1672)
);
defparam \d_cnst_sn.reg3_17_0[15] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[8]  (
	.I0(datai[8]),
	.I1(inf_abs0_2[8]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1665)
);
defparam \d_cnst_sn.reg3_17_0[8] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.un1_cf  (
	.I0(inf_abs0_2[23]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(\d_cnst_sn.reg3_5_sqmuxa_2_1 ),
	.I4(un87_df),
	.O(un1_cf)
);
defparam \d_cnst_sn.un1_cf .INIT=32'h04000000;
// @7:489
  LUT5 \d_cnst_sn.rd_4_sqmuxa  (
	.I0(inf_abs0_2[23]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un36_df),
	.I4(N_1890),
	.O(rd_4_sqmuxa)
);
defparam \d_cnst_sn.rd_4_sqmuxa .INIT=32'h00000001;
// @7:103
  LUT5 \d_cnst_sn.un1_df_16_2_RNISV2O2  (
	.I0(inf_abs0_2[23]),
	.I1(un1_b57),
	.I2(un1_df_17_2),
	.I3(un1_df_16),
	.I4(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.O(N_1841)
);
defparam \d_cnst_sn.un1_df_16_2_RNISV2O2 .INIT=32'h00BF0000;
// @7:103
  LUT4 \d_cnst_sn.un1_df_16  (
	.I0(inf_abs0_2[23]),
	.I1(un36_df),
	.I2(un1_b59),
	.I3(un87_df),
	.O(un1_df_16)
);
defparam \d_cnst_sn.un1_df_16 .INIT=16'h1000;
// @7:103
  LUT5 \d_cnst_sn.un1_b57_RNIEFGG1  (
	.I0(inf_abs0_2[23]),
	.I1(un1_b57),
	.I2(un36_df),
	.I3(un1_b59),
	.I4(un87_df),
	.O(N_1810)
);
defparam \d_cnst_sn.un1_b57_RNIEFGG1 .INIT=32'hFAFBFFFF;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_6_0_cZ[19]  (
	.I0(inf_abs0_2[28]),
	.I1(inf_abs0_2[29]),
	.I2(N_933),
	.I3(N_965),
	.I4(reg3_14_sqmuxa),
	.LO(\d_cnst_sn.reg3_17_6_0 [19])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[19] .INIT=32'hFD75FFFF;
// @7:103
  LUT3_L \d_cnst_sn.reg3_17_4_a2[13]  (
	.I0(inf_abs0_2[28]),
	.I1(reg3_14_sqmuxa),
	.I2(t_1[13]),
	.LO(reg3_17_4_a2[13])
);
defparam \d_cnst_sn.reg3_17_4_a2[13] .INIT=8'h40;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_3[2]  (
	.I0(inf_abs0_2[2]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[1]),
	.I3(reg3_14_sqmuxa),
	.I4(t_1[2]),
	.O(N_1752)
);
defparam \d_cnst_sn.reg3_17_3[2] .INIT=32'hC0AAF3AA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_3[1]  (
	.I0(inf_abs0_2[1]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[0]),
	.I3(reg3_14_sqmuxa),
	.I4(t_1[1]),
	.O(N_1751)
);
defparam \d_cnst_sn.reg3_17_3[1] .INIT=32'hC0AAF3AA;
// @7:103
  LUT4_L \d_cnst_sn.reg3_17_3[0]  (
	.I0(inf_abs0_2[0]),
	.I1(inf_abs0_2[28]),
	.I2(reg3_14_sqmuxa),
	.I3(t_1[0]),
	.LO(N_1750)
);
defparam \d_cnst_sn.reg3_17_3[0] .INIT=16'h0A3A;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_6_tz[24]  (
	.I0(inf_abs0_2[28]),
	.I1(r_4[23]),
	.I2(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I3(reg3_14_sqmuxa),
	.I4(N_1681),
	.O(\d_cnst_sn.reg3_17_0_tz [24])
);
defparam \d_cnst_sn.reg3_17_6_tz[24] .INIT=32'h8F0F8000;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_6_tz[22]  (
	.I0(inf_abs0_2[28]),
	.I1(r_4[21]),
	.I2(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I3(reg3_14_sqmuxa),
	.I4(N_1679),
	.O(\d_cnst_sn.reg3_17_0_tz [22])
);
defparam \d_cnst_sn.reg3_17_6_tz[22] .INIT=32'h8F0F8000;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_6_tz[23]  (
	.I0(inf_abs0_2[28]),
	.I1(r_4[22]),
	.I2(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I3(reg3_14_sqmuxa),
	.I4(N_1680),
	.O(\d_cnst_sn.reg3_17_0_tz [23])
);
defparam \d_cnst_sn.reg3_17_6_tz[23] .INIT=32'h8F0F8000;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_6_0_cZ[17]  (
	.I0(inf_abs0_2[17]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[16]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.LO(\d_cnst_sn.reg3_17_6_0 [17])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[17] .INIT=32'hF3F3AAFF;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_6_0_cZ[16]  (
	.I0(inf_abs0_2[16]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[15]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.LO(\d_cnst_sn.reg3_17_6_0 [16])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[16] .INIT=32'hF3F3AAFF;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_6_0_cZ[14]  (
	.I0(inf_abs0_2[14]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[13]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.LO(\d_cnst_sn.reg3_17_6_0 [14])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[14] .INIT=32'hF3F3AAFF;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_6_0_cZ[15]  (
	.I0(inf_abs0_2[15]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[14]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.LO(\d_cnst_sn.reg3_17_6_0 [15])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[15] .INIT=32'hF3F3AAFF;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_6_0_cZ[12]  (
	.I0(inf_abs0_2[12]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[11]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.LO(\d_cnst_sn.reg3_17_6_0 [12])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[12] .INIT=32'hF3F3AAFF;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_6_0_cZ[13]  (
	.I0(inf_abs0_2[13]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[12]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.LO(\d_cnst_sn.reg3_17_6_0 [13])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[13] .INIT=32'hF3F3AAFF;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_6_0_cZ[18]  (
	.I0(inf_abs0_2[18]),
	.I1(inf_abs0_2[28]),
	.I2(r_4[17]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.LO(\d_cnst_sn.reg3_17_6_0 [18])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[18] .INIT=32'hF3F3AAFF;
// @7:103
  LUT2 \d_cnst_sn.reg3_17_a1_2[21]  (
	.I0(inf_abs0_2[28]),
	.I1(reg3_14_sqmuxa),
	.O(\d_cnst_sn.reg3_17_a1_2 [24])
);
defparam \d_cnst_sn.reg3_17_a1_2[21] .INIT=4'h4;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[4]  (
	.I0(datai[4]),
	.I1(inf_abs0_2[4]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1661)
);
defparam \d_cnst_sn.reg3_17_0[4] .INIT=32'hAAACAAAA;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_0[3]  (
	.I0(datai[3]),
	.I1(inf_abs0_2[3]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.LO(N_1660)
);
defparam \d_cnst_sn.reg3_17_0[3] .INIT=32'hAAACAAAA;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_0[5]  (
	.I0(datai[5]),
	.I1(inf_abs0_2[5]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(un1_cf),
	.O(N_1662)
);
defparam \d_cnst_sn.reg3_17_0[5] .INIT=32'hAAACAAAA;
// @7:47
  LUT6 \d_cnst_sn.reg1_16_8_1837_3_1_cZ  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[26]),
	.I5(reg3_1_1[27]),
	.O(\d_cnst_sn.reg1_16_8_1837_3_1 )
);
defparam \d_cnst_sn.reg1_16_8_1837_3_1_cZ .INIT=64'hF8F8F0F808080008;
// @7:47
  LUT6 \d_cnst_sn.reg1_16_7_1870_3_1_cZ  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[25]),
	.I5(reg3_1_1[26]),
	.O(\d_cnst_sn.reg1_16_7_1870_3_1 )
);
defparam \d_cnst_sn.reg1_16_7_1870_3_1_cZ .INIT=64'hF8F8F0F808080008;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_9_2294_3_1_cZ  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[24]),
	.I5(reg3_1_1[25]),
	.O(\d_cnst_sn.reg0_28_9_2294_3_1 )
);
defparam \d_cnst_sn.reg0_28_9_2294_3_1_cZ .INIT=64'hF8F8F0F808080008;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_7_2360_3_1_cZ  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[22]),
	.I5(reg3_1_1[23]),
	.O(\d_cnst_sn.reg0_28_7_2360_3_1 )
);
defparam \d_cnst_sn.reg0_28_7_2360_3_1_cZ .INIT=64'hF8F8F0F808080008;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_6_2393_3_1_cZ  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[21]),
	.I5(reg3_1_1[22]),
	.O(\d_cnst_sn.reg0_28_6_2393_3_1 )
);
defparam \d_cnst_sn.reg0_28_6_2393_3_1_cZ .INIT=64'hF8F8F0F808080008;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_5_2426_3_1_cZ  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[20]),
	.I5(reg3_1_1[21]),
	.O(\d_cnst_sn.reg0_28_5_2426_3_1 )
);
defparam \d_cnst_sn.reg0_28_5_2426_3_1_cZ .INIT=64'hF8F8F0F808080008;
  LUT6 \d_cnst_sn.r_4_2_RNI0O8E1[18]  (
	.I0(reg0[18]),
	.I1(reg2[18]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_965),
	.O(r_4[18])
);
defparam \d_cnst_sn.r_4_2_RNI0O8E1[18] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNI0O8E1_0[18]  (
	.I0(reg0[18]),
	.I1(reg2[18]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_965),
	.O(un3_t_axb_18)
);
defparam \d_cnst_sn.r_4_2_RNI0O8E1_0[18] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIE8BE1_0[21]  (
	.I0(reg0[21]),
	.I1(reg2[21]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_968),
	.O(un3_t_axb_21)
);
defparam \d_cnst_sn.r_4_2_RNIE8BE1_0[21] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIE8BE1[21]  (
	.I0(reg0[21]),
	.I1(reg2[21]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_968),
	.O(r_4[21])
);
defparam \d_cnst_sn.r_4_2_RNIE8BE1[21] .INIT=64'hAFACAFAAA0ACA0AA;
// @7:358
  LUT5 un32_reg0_axb_29_cZ (
	.I0(datai[29]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[29]),
	.O(un32_reg0_axb_29)
);
defparam un32_reg0_axb_29_cZ.INIT=32'h2220DDDF;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_6[30]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[30]),
	.I5(reg3_1_1[30]),
	.O(N_1493)
);
defparam \d_cnst_sn.reg2_16_6[30] .INIT=64'hFF0DFF01000C0000;
// @7:74
  LUT6 \d_cnst_sn.reg2_16[28]  (
	.I0(un3_reg3_s_25),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[28]),
	.I5(reg3_1_1[28]),
	.O(N_1363)
);
defparam \d_cnst_sn.reg2_16[28] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16[27]  (
	.I0(un3_reg3_s_24),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[27]),
	.I5(reg3_1_1[27]),
	.O(N_1362)
);
defparam \d_cnst_sn.reg2_16[27] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16[26]  (
	.I0(un3_reg3_s_23),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[26]),
	.I5(reg3_1_1[26]),
	.O(N_1361)
);
defparam \d_cnst_sn.reg2_16[26] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[19]  (
	.I0(un3_reg3_s_16),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[19]),
	.I5(reg3_1_1[19]),
	.O(N_1354)
);
defparam \d_cnst_sn.reg2_16_2[19] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[18]  (
	.I0(un3_reg3_s_15),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[18]),
	.I5(reg3_1_1[18]),
	.O(N_1353)
);
defparam \d_cnst_sn.reg2_16_2[18] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[17]  (
	.I0(un3_reg3_s_14),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[17]),
	.I5(reg3_1_1[17]),
	.O(N_1352)
);
defparam \d_cnst_sn.reg2_16_2[17] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[16]  (
	.I0(un3_reg3_s_13),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[16]),
	.I5(reg3_1_1[16]),
	.O(N_1351)
);
defparam \d_cnst_sn.reg2_16_2[16] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[15]  (
	.I0(un3_reg3_s_12),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[15]),
	.I5(reg3_1_1[15]),
	.O(N_1350)
);
defparam \d_cnst_sn.reg2_16_2[15] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[14]  (
	.I0(un3_reg3_s_11),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[14]),
	.I5(reg3_1_1[14]),
	.O(N_1349)
);
defparam \d_cnst_sn.reg2_16_2[14] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[13]  (
	.I0(un3_reg3_s_10),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[13]),
	.I5(reg3_1_1[13]),
	.O(N_1348)
);
defparam \d_cnst_sn.reg2_16_2[13] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[12]  (
	.I0(un3_reg3_s_9),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[12]),
	.I5(reg3_1_1[12]),
	.O(N_1347)
);
defparam \d_cnst_sn.reg2_16_2[12] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[11]  (
	.I0(un3_reg3_s_8),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[11]),
	.I5(reg3_1_1[11]),
	.O(N_1346)
);
defparam \d_cnst_sn.reg2_16_2[11] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[10]  (
	.I0(un3_reg3_s_7),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[10]),
	.I5(reg3_1_1[10]),
	.O(N_1345)
);
defparam \d_cnst_sn.reg2_16_2[10] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[9]  (
	.I0(un3_reg3_s_6),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[9]),
	.I5(reg3_1_1[9]),
	.O(N_1344)
);
defparam \d_cnst_sn.reg2_16_2[9] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[8]  (
	.I0(un3_reg3_s_5),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[8]),
	.I5(reg3_1_1[8]),
	.O(N_1343)
);
defparam \d_cnst_sn.reg2_16_2[8] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[7]  (
	.I0(un3_reg3_s_4),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[7]),
	.I5(reg3_1_1[7]),
	.O(N_1342)
);
defparam \d_cnst_sn.reg2_16_2[7] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[6]  (
	.I0(un3_reg3_s_3),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[6]),
	.I5(reg3_1_1[6]),
	.O(N_1341)
);
defparam \d_cnst_sn.reg2_16_2[6] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[5]  (
	.I0(un3_reg3_s_2),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[5]),
	.I5(reg3_1_1[5]),
	.O(N_1340)
);
defparam \d_cnst_sn.reg2_16_2[5] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[4]  (
	.I0(un3_reg3_s_1),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[4]),
	.I5(reg3_1_1[4]),
	.O(N_1339)
);
defparam \d_cnst_sn.reg2_16_2[4] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[3]  (
	.I0(reg3[3]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[3]),
	.I5(reg3_1_1[3]),
	.O(N_1338)
);
defparam \d_cnst_sn.reg2_16_2[3] .INIT=64'hFFF7FF0700F40004;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[2]  (
	.I0(reg3[2]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[2]),
	.I5(reg3_1_1[2]),
	.O(N_1337)
);
defparam \d_cnst_sn.reg2_16_2[2] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2[1]  (
	.I0(reg3[1]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[1]),
	.I5(reg3_1_1[1]),
	.O(N_1336)
);
defparam \d_cnst_sn.reg2_16_2[1] .INIT=64'hFFFBFF0B00F80008;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_1_0[25]  (
	.I0(un3_reg3_s_22),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[31]),
	.I3(\d_cnst_sn.reg0_28_a0_1 [7]),
	.I4(\d_cnst_sn.reg2_16_0 [25]),
	.I5(reg3_1_1[25]),
	.O(\d_cnst_sn.reg2_16_1 [25])
);
defparam \d_cnst_sn.reg2_16_1_0[25] .INIT=64'hFBFF000008FF0000;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_1_0[24]  (
	.I0(un3_reg3_s_21),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[31]),
	.I3(\d_cnst_sn.reg0_28_a0_1 [7]),
	.I4(\d_cnst_sn.reg2_16_0 [24]),
	.I5(reg3_1_1[24]),
	.O(\d_cnst_sn.reg2_16_1 [24])
);
defparam \d_cnst_sn.reg2_16_1_0[24] .INIT=64'hFBFF000008FF0000;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_1_0[23]  (
	.I0(un3_reg3_s_20),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[31]),
	.I3(\d_cnst_sn.reg0_28_a0_1 [7]),
	.I4(\d_cnst_sn.reg2_16_0 [23]),
	.I5(reg3_1_1[23]),
	.O(\d_cnst_sn.reg2_16_1 [23])
);
defparam \d_cnst_sn.reg2_16_1_0[23] .INIT=64'hFBFF000008FF0000;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_1_0[22]  (
	.I0(un3_reg3_s_19),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[31]),
	.I3(\d_cnst_sn.reg0_28_a0_1 [7]),
	.I4(\d_cnst_sn.reg2_16_0 [22]),
	.I5(reg3_1_1[22]),
	.O(\d_cnst_sn.reg2_16_1 [22])
);
defparam \d_cnst_sn.reg2_16_1_0[22] .INIT=64'hFBFF000008FF0000;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_1_0[21]  (
	.I0(un3_reg3_s_18),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[31]),
	.I3(\d_cnst_sn.reg0_28_a0_1 [7]),
	.I4(reg3_1_1[21]),
	.I5(\d_cnst_sn.reg2_16_0 [21]),
	.O(\d_cnst_sn.reg2_16_1 [21])
);
defparam \d_cnst_sn.reg2_16_1_0[21] .INIT=64'hFBFF08FF00000000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_0[16]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[15]),
	.I4(reg3_1_1[16]),
	.I5(t_1[16]),
	.O(N_1083)
);
defparam \d_cnst_sn.reg0_28_0[16] .INIT=64'hFDDD2000FFDF2202;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_0[15]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[14]),
	.I4(reg3_1_1[15]),
	.I5(t_1[15]),
	.O(N_1082)
);
defparam \d_cnst_sn.reg0_28_0[15] .INIT=64'hFDDD2000FFDF2202;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_0[14]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[13]),
	.I4(reg3_1_1[14]),
	.I5(t_1[14]),
	.O(N_1081)
);
defparam \d_cnst_sn.reg0_28_0[14] .INIT=64'hFDDD2000FFDF2202;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_0[13]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[12]),
	.I4(reg3_1_1[13]),
	.I5(t_1[13]),
	.O(N_1080)
);
defparam \d_cnst_sn.reg0_28_0[13] .INIT=64'hFDDD2000FFDF2202;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_0[12]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[11]),
	.I4(reg3_1_1[12]),
	.I5(t_1[12]),
	.O(N_1079)
);
defparam \d_cnst_sn.reg0_28_0[12] .INIT=64'hFDDD2000FFDF2202;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_0[11]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[10]),
	.I4(reg3_1_1[11]),
	.I5(t_1[11]),
	.O(N_1078)
);
defparam \d_cnst_sn.reg0_28_0[11] .INIT=64'hFDDD2000FFDF2202;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_0[10]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[9]),
	.I4(reg3_1_1[10]),
	.I5(t_1[10]),
	.O(N_1077)
);
defparam \d_cnst_sn.reg0_28_0[10] .INIT=64'hFDDD2000FFDF2202;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_0[9]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[8]),
	.I4(reg3_1_1[9]),
	.I5(t_1[9]),
	.O(N_1076)
);
defparam \d_cnst_sn.reg0_28_0[9] .INIT=64'hFDDD2000FFDF2202;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_7[2]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(reg3_1_1[2]),
	.I4(r_4[1]),
	.I5(t_1[2]),
	.LO(N_1069)
);
defparam \d_cnst_sn.reg0_28_7[2] .INIT=64'hFD20DD00FF22DF02;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_7[1]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(reg3_1_1[1]),
	.I4(r_4[0]),
	.I5(t_1[1]),
	.O(N_1068)
);
defparam \d_cnst_sn.reg0_28_7[1] .INIT=64'hFD20DD00FF22DF02;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_14_0_cZ  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(N_3568),
	.I5(reg3_1_1[30]),
	.O(\d_cnst_sn.reg0_28_14_0 )
);
defparam \d_cnst_sn.reg0_28_14_0_cZ .INIT=64'hFFFFC101FFFF0000;
  LUT6 \d_cnst_sn.r_4_RNITKAH1[4]  (
	.I0(reg1[4]),
	.I1(un3_reg3_s_1),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_919),
	.O(r_4[4])
);
defparam \d_cnst_sn.r_4_RNITKAH1[4] .INIT=64'hFCFFFAFF0C000A00;
  LUT6 \d_cnst_sn.r_4_RNITKAH1_0[4]  (
	.I0(reg1[4]),
	.I1(un3_reg3_s_1),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_919),
	.O(un3_t_axb_4)
);
defparam \d_cnst_sn.r_4_RNITKAH1_0[4] .INIT=64'h03000500F3FFF5FF;
  LUT6 \d_cnst_sn.r_4_RNI9T9D1_0[1]  (
	.I0(reg1[1]),
	.I1(reg3[1]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_916),
	.O(un3_t_axb_1)
);
defparam \d_cnst_sn.r_4_RNI9T9D1_0[1] .INIT=64'h03000500F3FFF5FF;
  LUT6 \d_cnst_sn.r_4_RNI9T9D1[1]  (
	.I0(reg1[1]),
	.I1(reg3[1]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_916),
	.O(r_4[1])
);
defparam \d_cnst_sn.r_4_RNI9T9D1[1] .INIT=64'hFCFFFAFF0C000A00;
  LUT6 \d_cnst_sn.r_4_RNI6Q9D1[0]  (
	.I0(reg1[0]),
	.I1(reg3[0]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_915),
	.O(r_4[0])
);
defparam \d_cnst_sn.r_4_RNI6Q9D1[0] .INIT=64'hFCFFFAFF0C000A00;
  LUT6 \d_cnst_sn.r_4_RNI6Q9D1_0[0]  (
	.I0(reg1[0]),
	.I1(reg3[0]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_915),
	.O(un3_t_axb_0)
);
defparam \d_cnst_sn.r_4_RNI6Q9D1_0[0] .INIT=64'h03000500F3FFF5FF;
  LUT6 \d_cnst_sn.r_4_1_RNI3T3N1[24]  (
	.I0(reg1[24]),
	.I1(un3_reg3_s_21),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_939),
	.O(r_4[24])
);
defparam \d_cnst_sn.r_4_1_RNI3T3N1[24] .INIT=64'hFCFFFAFF0C000A00;
  LUT6 \d_cnst_sn.r_4_1_RNI3T3N1_0[24]  (
	.I0(reg1[24]),
	.I1(un3_reg3_s_21),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_939),
	.O(un3_t_axb_24)
);
defparam \d_cnst_sn.r_4_1_RNI3T3N1_0[24] .INIT=64'h03000500F3FFF5FF;
  LUT6 \d_cnst_sn.r_4_1_RNI0R3N1[23]  (
	.I0(reg1[23]),
	.I1(un3_reg3_s_20),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_938),
	.O(r_4[23])
);
defparam \d_cnst_sn.r_4_1_RNI0R3N1[23] .INIT=64'hFCFFFAFF0C000A00;
  LUT6 \d_cnst_sn.r_4_1_RNI0R3N1_0[23]  (
	.I0(reg1[23]),
	.I1(un3_reg3_s_20),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_938),
	.O(un3_t_axb_23)
);
defparam \d_cnst_sn.r_4_1_RNI0R3N1_0[23] .INIT=64'h03000500F3FFF5FF;
  LUT6 \d_cnst_sn.r_4_1_RNIC34N1[27]  (
	.I0(reg1[27]),
	.I1(un3_reg3_s_24),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_942),
	.O(r_4[27])
);
defparam \d_cnst_sn.r_4_1_RNIC34N1[27] .INIT=64'hFCFFFAFF0C000A00;
  LUT6 \d_cnst_sn.r_4_1_RNIC34N1_0[27]  (
	.I0(reg1[27]),
	.I1(un3_reg3_s_24),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_942),
	.O(un3_t_axb_27)
);
defparam \d_cnst_sn.r_4_1_RNIC34N1_0[27] .INIT=64'h03000500F3FFF5FF;
  LUT6 \d_cnst_sn.r_4_1_RNI0K3N1[20]  (
	.I0(reg1[20]),
	.I1(un3_reg3_s_17),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_935),
	.O(r_4[20])
);
defparam \d_cnst_sn.r_4_1_RNI0K3N1[20] .INIT=64'hFCFFFAFF0C000A00;
  LUT6 \d_cnst_sn.r_4_1_RNI0K3N1_0[20]  (
	.I0(reg1[20]),
	.I1(un3_reg3_s_17),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_935),
	.O(un3_t_axb_20)
);
defparam \d_cnst_sn.r_4_1_RNI0K3N1_0[20] .INIT=64'h03000500F3FFF5FF;
  LUT6 \d_cnst_sn.r_4_2_RNIQKBE1[25]  (
	.I0(reg0[25]),
	.I1(reg2[25]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_972),
	.O(r_4[25])
);
defparam \d_cnst_sn.r_4_2_RNIQKBE1[25] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNIQKBE1_0[25]  (
	.I0(reg0[25]),
	.I1(reg2[25]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_972),
	.O(un3_t_axb_25)
);
defparam \d_cnst_sn.r_4_2_RNIQKBE1_0[25] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNI3UBE1[28]  (
	.I0(reg0[28]),
	.I1(reg2[28]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_975),
	.O(r_4[28])
);
defparam \d_cnst_sn.r_4_2_RNI3UBE1[28] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNI3UBE1_0[28]  (
	.I0(reg0[28]),
	.I1(reg2[28]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_975),
	.O(un3_t_axb_28)
);
defparam \d_cnst_sn.r_4_2_RNI3UBE1_0[28] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNITNBE1[26]  (
	.I0(reg0[26]),
	.I1(reg2[26]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_973),
	.O(r_4[26])
);
defparam \d_cnst_sn.r_4_2_RNITNBE1[26] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNITNBE1_0[26]  (
	.I0(reg0[26]),
	.I1(reg2[26]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_973),
	.O(un3_t_axb_26)
);
defparam \d_cnst_sn.r_4_2_RNITNBE1_0[26] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_1_RNI6O3N1_0[22]  (
	.I0(reg1[22]),
	.I1(un3_reg3_s_19),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_937),
	.O(un3_t_axb_22)
);
defparam \d_cnst_sn.r_4_1_RNI6O3N1_0[22] .INIT=64'h03000500F3FFF5FF;
  LUT6 \d_cnst_sn.r_4_1_RNI6O3N1[22]  (
	.I0(reg1[22]),
	.I1(un3_reg3_s_19),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_937),
	.O(r_4[22])
);
defparam \d_cnst_sn.r_4_1_RNI6O3N1[22] .INIT=64'hFCFFFAFF0C000A00;
  LUT6 \d_cnst_sn.r_4_RNIF3AD1[3]  (
	.I0(reg1[3]),
	.I1(reg3[3]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_918),
	.O(r_4[3])
);
defparam \d_cnst_sn.r_4_RNIF3AD1[3] .INIT=64'hF3FFFAFF03000A00;
  LUT6 \d_cnst_sn.r_4_RNIF3AD1_0[3]  (
	.I0(reg1[3]),
	.I1(reg3[3]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_918),
	.O(un3_t_axb_3)
);
defparam \d_cnst_sn.r_4_RNIF3AD1_0[3] .INIT=64'h0C000500FCFFF5FF;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_a2_2_0_cZ[21]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_967),
	.I4(N_935),
	.O(\d_cnst_sn.reg3_17_a2_2_0 [21])
);
defparam \d_cnst_sn.reg3_17_a2_2_0_cZ[21] .INIT=32'h44044000;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_4_a2_0_cZ[27]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_941),
	.I4(N_973),
	.O(\d_cnst_sn.reg3_17_4_a2_0 [27])
);
defparam \d_cnst_sn.reg3_17_4_a2_0_cZ[27] .INIT=32'h44400400;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_4_a2_0_cZ[25]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_971),
	.I4(N_939),
	.O(\d_cnst_sn.reg3_17_4_a2_0 [25])
);
defparam \d_cnst_sn.reg3_17_4_a2_0_cZ[25] .INIT=32'h44044000;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_4_a2_0_cZ[28]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_974),
	.I4(N_942),
	.O(\d_cnst_sn.reg3_17_4_a2_0 [28])
);
defparam \d_cnst_sn.reg3_17_4_a2_0_cZ[28] .INIT=32'h44044000;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_4_a2_0_cZ[26]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_940),
	.I4(N_972),
	.O(\d_cnst_sn.reg3_17_4_a2_0 [26])
);
defparam \d_cnst_sn.reg3_17_4_a2_0_cZ[26] .INIT=32'h44400400;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_7_d[24]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_970),
	.I4(N_938),
	.I5(reg3_1_1[24]),
	.O(reg0_28_7_d[24])
);
defparam \d_cnst_sn.reg0_28_7_d[24] .INIT=64'hFFDFFDDD22022000;
  LUT6 \datai_RNIL2NH1[26]  (
	.I0(datai[26]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_941),
	.I4(N_973),
	.I5(m7),
	.O(un32_reg0_axb_26)
);
defparam \datai_RNIL2NH1[26] .INIT=64'h00CF30FFAA659A55;
  LUT6 \datai_RNIIVMH1[25]  (
	.I0(datai[25]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_940),
	.I4(N_972),
	.I5(m7),
	.O(un32_reg0_axb_25)
);
defparam \datai_RNIIVMH1[25] .INIT=64'h00CF30FFAA659A55;
  LUT6 \d_cnst_sn.r_4_2_RNICPMH1[23]  (
	.I0(datai[23]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_970),
	.I4(N_938),
	.I5(m7),
	.O(un32_reg0_axb_23)
);
defparam \d_cnst_sn.r_4_2_RNICPMH1[23] .INIT=64'h0030CFFFAA9A6555;
  LUT6 \d_cnst_sn.r_4_0_0_RNID9G41[1]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(r_4_2_a0[1]),
	.I3(\d_cnst_sn.r_4_0_0 [1]),
	.I4(N_916),
	.I5(m_2[1]),
	.O(un32_reg0_axb_1)
);
defparam \d_cnst_sn.r_4_0_0_RNID9G41[1] .INIT=64'hBFBB04004044FBFF;
  LUT6 \d_cnst_sn.r_4_2_a0_RNI4HHP2[0]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(m_2_i[0]),
	.I3(r_4_2_a0[0]),
	.I4(\d_cnst_sn.r_4_0_0 [0]),
	.I5(N_915),
	.O(N_1035)
);
defparam \d_cnst_sn.r_4_2_a0_RNI4HHP2[0] .INIT=64'h4B0F4B4BF0B4F0F0;
  LUT6 \datai_RNIR8NH1[28]  (
	.I0(datai[28]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_943),
	.I4(N_975),
	.I5(m7),
	.O(un32_reg0_axb_28)
);
defparam \datai_RNIR8NH1[28] .INIT=64'h00CF30FFAA659A55;
  LUT6 \d_cnst_sn.r_4_2_RNIO5NH1[27]  (
	.I0(datai[27]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_974),
	.I4(N_942),
	.I5(m7),
	.O(un32_reg0_axb_27)
);
defparam \d_cnst_sn.r_4_2_RNIO5NH1[27] .INIT=64'h0030CFFFAA9A6555;
  LUT6 \datai_RNI3GMH1[20]  (
	.I0(datai[20]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_967),
	.I4(N_935),
	.I5(m7),
	.O(un32_reg0_axb_20)
);
defparam \datai_RNI3GMH1[20] .INIT=64'h0030CFFFAA9A6555;
  LUT6 \d_cnst_sn.r_4_2_RNIFSMH1[24]  (
	.I0(datai[24]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_971),
	.I4(N_939),
	.I5(m7),
	.O(un32_reg0_axb_24)
);
defparam \d_cnst_sn.r_4_2_RNIFSMH1[24] .INIT=64'h0030CFFFAA9A6555;
  LUT6 \datai_RNI9MMH1[22]  (
	.I0(datai[22]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_969),
	.I4(N_937),
	.I5(m7),
	.O(un32_reg0_axb_22)
);
defparam \datai_RNI9MMH1[22] .INIT=64'h0030CFFFAA9A6555;
  LUT6 \d_cnst_sn.r_4_1_RNI6JMH1[21]  (
	.I0(datai[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[29]),
	.I3(N_936),
	.I4(N_968),
	.I5(m7),
	.O(un32_reg0_axb_21)
);
defparam \d_cnst_sn.r_4_1_RNI6JMH1[21] .INIT=64'h00CF30FFAA659A55;
// @7:47
  LUT5 \dce_cZ[0]  (
	.I0(state[0]),
	.I1(inf_abs0_2[23]),
	.I2(inf_abs0_2[31]),
	.I3(un1_df_1),
	.I4(un36_df),
	.O(dce[0])
);
defparam \dce_cZ[0] .INIT=32'h000000A2;
// @7:74
  LUT6 \d_cnst_sn.un1_state_4_1  (
	.I0(state[0]),
	.I1(inf_abs0_2[23]),
	.I2(inf_abs0_2[31]),
	.I3(N_1892),
	.I4(un36_df),
	.I5(N_1890),
	.O(\d_cnst_sn.un1_state_3_1 )
);
defparam \d_cnst_sn.un1_state_4_1 .INIT=64'hFFFFFF5DFFFFFFFF;
// @7:103
  LUT4 \d_cnst_sn.reg3_m2_7  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(N_28),
	.I3(t_1[3]),
	.O(t_6[3])
);
defparam \d_cnst_sn.reg3_m2_7 .INIT=16'h40FB;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_12_2195_a6  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(N_1033),
	.I4(un32_reg0_s_28),
	.I5(un11_reg0_s_28),
	.O(N_3614)
);
defparam \d_cnst_sn.reg0_28_12_2195_a6 .INIT=64'h0606060000060000;
// @7:318
  LUT5 un11_reg0_axb_29_cZ (
	.I0(datai[29]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[29]),
	.O(un11_reg0_axb_29)
);
defparam un11_reg0_axb_29_cZ.INIT=32'hDDDF2220;
  LUT6 \d_cnst_sn.r_4_3[19]  (
	.I0(reg0[19]),
	.I1(reg2[19]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_2722),
	.O(r_4[19])
);
defparam \d_cnst_sn.r_4_3[19] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_3_i[19]  (
	.I0(reg0[19]),
	.I1(reg2[19]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_2722),
	.O(un3_t_axb_19)
);
defparam \d_cnst_sn.r_4_3_i[19] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNI7PRB1[6]  (
	.I0(reg0[6]),
	.I1(reg2[6]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_953),
	.O(r_4[6])
);
defparam \d_cnst_sn.r_4_2_RNI7PRB1[6] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNI7PRB1_0[6]  (
	.I0(reg0[6]),
	.I1(reg2[6]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_953),
	.O(un3_t_axb_6)
);
defparam \d_cnst_sn.r_4_2_RNI7PRB1_0[6] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIE58E1_0[12]  (
	.I0(reg0[12]),
	.I1(reg2[12]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_959),
	.O(un3_t_axb_12)
);
defparam \d_cnst_sn.r_4_2_RNIE58E1_0[12] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIE58E1[12]  (
	.I0(reg0[12]),
	.I1(reg2[12]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_959),
	.O(r_4[12])
);
defparam \d_cnst_sn.r_4_2_RNIE58E1[12] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNI4MRB1[5]  (
	.I0(reg0[5]),
	.I1(reg2[5]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_952),
	.O(r_4[5])
);
defparam \d_cnst_sn.r_4_2_RNI4MRB1[5] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNI4MRB1_0[5]  (
	.I0(reg0[5]),
	.I1(reg2[5]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_952),
	.O(un3_t_axb_5)
);
defparam \d_cnst_sn.r_4_2_RNI4MRB1_0[5] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNITK8E1[17]  (
	.I0(reg0[17]),
	.I1(reg2[17]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_964),
	.O(r_4[17])
);
defparam \d_cnst_sn.r_4_2_RNITK8E1[17] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNITK8E1_0[17]  (
	.I0(reg0[17]),
	.I1(reg2[17]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_964),
	.O(un3_t_axb_17)
);
defparam \d_cnst_sn.r_4_2_RNITK8E1_0[17] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIASRB1[7]  (
	.I0(reg0[7]),
	.I1(reg2[7]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_954),
	.O(r_4[7])
);
defparam \d_cnst_sn.r_4_2_RNIASRB1[7] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNIASRB1_0[7]  (
	.I0(reg0[7]),
	.I1(reg2[7]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_954),
	.O(un3_t_axb_7)
);
defparam \d_cnst_sn.r_4_2_RNIASRB1_0[7] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIG2SB1[9]  (
	.I0(reg0[9]),
	.I1(reg2[9]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_956),
	.O(r_4[9])
);
defparam \d_cnst_sn.r_4_2_RNIG2SB1[9] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNIG2SB1_0[9]  (
	.I0(reg0[9]),
	.I1(reg2[9]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_956),
	.O(un3_t_axb_9)
);
defparam \d_cnst_sn.r_4_2_RNIG2SB1_0[9] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNI8V7E1[10]  (
	.I0(reg0[10]),
	.I1(reg2[10]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_957),
	.O(r_4[10])
);
defparam \d_cnst_sn.r_4_2_RNI8V7E1[10] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNI8V7E1_0[10]  (
	.I0(reg0[10]),
	.I1(reg2[10]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_957),
	.O(un3_t_axb_10)
);
defparam \d_cnst_sn.r_4_2_RNI8V7E1_0[10] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIKB8E1_0[14]  (
	.I0(reg0[14]),
	.I1(reg2[14]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_961),
	.O(un3_t_axb_14)
);
defparam \d_cnst_sn.r_4_2_RNIKB8E1_0[14] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIKB8E1[14]  (
	.I0(reg0[14]),
	.I1(reg2[14]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_961),
	.O(r_4[14])
);
defparam \d_cnst_sn.r_4_2_RNIKB8E1[14] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNIQH8E1[16]  (
	.I0(reg0[16]),
	.I1(reg2[16]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_963),
	.O(r_4[16])
);
defparam \d_cnst_sn.r_4_2_RNIQH8E1[16] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNIQH8E1_0[16]  (
	.I0(reg0[16]),
	.I1(reg2[16]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_963),
	.O(un3_t_axb_16)
);
defparam \d_cnst_sn.r_4_2_RNIQH8E1_0[16] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIH88E1[13]  (
	.I0(reg0[13]),
	.I1(reg2[13]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_960),
	.O(r_4[13])
);
defparam \d_cnst_sn.r_4_2_RNIH88E1[13] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNIH88E1_0[13]  (
	.I0(reg0[13]),
	.I1(reg2[13]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_960),
	.O(un3_t_axb_13)
);
defparam \d_cnst_sn.r_4_2_RNIH88E1_0[13] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_2_RNIB28E1[11]  (
	.I0(reg0[11]),
	.I1(reg2[11]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_958),
	.O(r_4[11])
);
defparam \d_cnst_sn.r_4_2_RNIB28E1[11] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNIB28E1_0[11]  (
	.I0(reg0[11]),
	.I1(reg2[11]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_958),
	.O(un3_t_axb_11)
);
defparam \d_cnst_sn.r_4_2_RNIB28E1_0[11] .INIT=64'h505350555F535F55;
  LUT6 \d_cnst_sn.r_4_0_0_0_RNIFROS1[4]  (
	.I0(reg1[4]),
	.I1(inf_abs0_2[30]),
	.I2(\d_cnst_sn.r_4_0_0 [4]),
	.I3(N_919),
	.I4(m_2[4]),
	.I5(N_13),
	.O(un32_reg0_axb_4)
);
defparam \d_cnst_sn.r_4_0_0_0_RNIFROS1[4] .INIT=64'hFF0000FFE0E01F1F;
  LUT6 \d_cnst_sn.r_4_2_RNINE8E1[15]  (
	.I0(reg0[15]),
	.I1(reg2[15]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_962),
	.O(r_4[15])
);
defparam \d_cnst_sn.r_4_2_RNINE8E1[15] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNINE8E1_0[15]  (
	.I0(reg0[15]),
	.I1(reg2[15]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_962),
	.O(un3_t_axb_15)
);
defparam \d_cnst_sn.r_4_2_RNINE8E1_0[15] .INIT=64'h505350555F535F55;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_8_627_i_1_RNIKNJN1  (
	.I0(state[0]),
	.I1(un1_inf_abs0_10[1]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(\d_cnst_sn.addr_20_iv_8_627_i_1 ),
	.I5(N_2641),
	.LO(N_2315_i)
);
defparam \d_cnst_sn.addr_20_iv_8_627_i_1_RNIKNJN1 .INIT=64'h000000000000DFFF;
  LUT6 \d_cnst_sn.r_4_2_RNIDVRB1[8]  (
	.I0(reg0[8]),
	.I1(reg2[8]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_955),
	.O(r_4[8])
);
defparam \d_cnst_sn.r_4_2_RNIDVRB1[8] .INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 \d_cnst_sn.r_4_2_RNIDVRB1_0[8]  (
	.I0(reg0[8]),
	.I1(reg2[8]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.I5(N_955),
	.O(un3_t_axb_8)
);
defparam \d_cnst_sn.r_4_2_RNIDVRB1_0[8] .INIT=64'h505350555F535F55;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_7_654_i_1_RNIG3SC1  (
	.I0(reg2[0]),
	.I1(inf_abs0_2[0]),
	.I2(inf_abs0_2[28]),
	.I3(\d_cnst_sn.addr_20_iv_7_654_i_1 ),
	.I4(N_2660_2),
	.I5(N_2641),
	.LO(N_2335_i)
);
defparam \d_cnst_sn.addr_20_iv_7_654_i_1_RNIG3SC1 .INIT=64'h00000000006F00FF;
  LUT6 \d_cnst_sn.r_4_0_0_0_RNIBNOS1[3]  (
	.I0(reg1[3]),
	.I1(inf_abs0_2[30]),
	.I2(\d_cnst_sn.r_4_0_0 [3]),
	.I3(N_918),
	.I4(m_2[3]),
	.I5(N_13),
	.O(un32_reg0_axb_3)
);
defparam \d_cnst_sn.r_4_0_0_0_RNIBNOS1[3] .INIT=64'hFF0000FFE0E01F1F;
  LUT6 \datai_RNIO9B94[2]  (
	.I0(datai[2]),
	.I1(inf_abs0_2[2]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(N_28),
	.O(un32_reg0_axb_2)
);
defparam \datai_RNIO9B94[2] .INIT=64'hCACACACC35353533;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[22]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_22),
	.I3(un11_reg0_s_22),
	.O(N_1581)
);
defparam \d_cnst_sn.reg2_16_9[22] .INIT=16'hFD20;
// @7:118
  LUT6 un11_r_df22_cZ (
	.I0(N_969),
	.I1(N_937),
	.I2(m_2[22]),
	.I3(m_2[23]),
	.I4(N_13),
	.I5(r_4[23]),
	.O(un11_r_df22)
);
defparam un11_r_df22_cZ.INIT=64'hC300A50000C300A5;
// @7:118
  LUT6 un11_r_lt22_cZ (
	.I0(N_969),
	.I1(N_937),
	.I2(m_2[22]),
	.I3(m_2[23]),
	.I4(N_13),
	.I5(r_4[23]),
	.O(un11_r_lt22)
);
defparam un11_r_lt22_cZ.INIT=64'h30005000FF30FF50;
// @7:151
  LUT6 un26_r_lt22_cZ (
	.I0(N_969),
	.I1(N_937),
	.I2(m_2[22]),
	.I3(m_2[23]),
	.I4(N_13),
	.I5(r_4[23]),
	.O(un26_r_lt22)
);
defparam un26_r_lt22_cZ.INIT=64'h30005000FF30FF50;
// @7:151
  LUT6 un26_r_df22_cZ (
	.I0(N_969),
	.I1(N_937),
	.I2(m_2[22]),
	.I3(m_2[23]),
	.I4(N_13),
	.I5(r_4[23]),
	.O(un26_r_df22)
);
defparam un26_r_df22_cZ.INIT=64'hC300A50000C300A5;
// @7:143
  LUT6 b18_df22_cZ (
	.I0(N_969),
	.I1(N_937),
	.I2(m_2[22]),
	.I3(m_2[23]),
	.I4(N_13),
	.I5(r_4[23]),
	.O(b18_df22)
);
defparam b18_df22_cZ.INIT=64'hC300A50000C300A5;
// @7:143
  LUT6 b18_lt22_cZ (
	.I0(N_969),
	.I1(N_937),
	.I2(m_2[22]),
	.I3(m_2[23]),
	.I4(N_13),
	.I5(r_4[23]),
	.O(b18_lt22)
);
defparam b18_lt22_cZ.INIT=64'h0CFF0AFF000C000A;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[8]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_8),
	.I3(un11_reg0_s_8),
	.O(N_1375)
);
defparam \d_cnst_sn.reg2_16_3[8] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[23]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_23),
	.I3(un11_reg0_s_23),
	.O(N_1582)
);
defparam \d_cnst_sn.reg2_16_9[23] .INIT=16'hFD20;
// @7:103
  LUT4_L \d_cnst_sn.b_cnst_0_m2_0  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(b18),
	.I3(un26_r_cry[30]),
	.LO(N_895)
);
defparam \d_cnst_sn.b_cnst_0_m2_0 .INIT=16'h2F0D;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[21]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_21),
	.I3(un11_reg0_s_21),
	.O(N_1580)
);
defparam \d_cnst_sn.reg2_16_9[21] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[16]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_16),
	.I3(un11_reg0_s_16),
	.O(N_1575)
);
defparam \d_cnst_sn.reg2_16_9[16] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[14]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_14),
	.I3(un11_reg0_s_14),
	.O(N_1381)
);
defparam \d_cnst_sn.reg2_16_3[14] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[24]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_24),
	.I3(un11_reg0_s_24),
	.O(N_1583)
);
defparam \d_cnst_sn.reg2_16_9[24] .INIT=16'hFD20;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[2]  (
	.I0(r_4_2_a0[1]),
	.I1(\d_cnst_sn.r_4_0_0 [1]),
	.I2(N_916),
	.I3(N_527_i),
	.I4(N_13),
	.I5(t_1[2]),
	.LO(t_6[2])
);
defparam \d_cnst_sn.reg2_16_11_RNO[2] .INIT=64'hF0004400F0FF44FF;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[2]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un11_reg0_s_2),
	.I3(un32_reg0_s_2),
	.O(N_1369)
);
defparam \d_cnst_sn.reg2_16_3[2] .INIT=16'hF2D0;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[5]  (
	.I0(r_4_2_a1_lut6_2_O5[3]),
	.I1(\d_cnst_sn.r_4_0_0 [4]),
	.I2(N_919),
	.I3(N_527_i),
	.I4(N_13),
	.I5(t_1[5]),
	.LO(t_6[5])
);
defparam \d_cnst_sn.reg2_16_11_RNO[5] .INIT=64'hF0004400F0FF44FF;
// @7:103
  LUT6_L \d_cnst_sn.r_4_2_a1_lut6_2_RNI5V8R3[3]  (
	.I0(r_4_2_a1_lut6_2_O5[3]),
	.I1(\d_cnst_sn.r_4_0_0 [4]),
	.I2(N_919),
	.I3(N_527_i),
	.I4(N_13),
	.I5(t_1[5]),
	.LO(r_4_2_a1_lut6_2_RNI5V8R3[3])
);
defparam \d_cnst_sn.r_4_2_a1_lut6_2_RNI5V8R3[3] .INIT=64'h0FFFBBFF0F00BB00;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_21_1130_i_m2  (
	.I0(reg1[19]),
	.I1(reg0[19]),
	.I2(reg2[19]),
	.I3(un3_reg3_s_16),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(N_2724)
);
defparam \d_cnst_sn.r_4_3_21_1130_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[4]  (
	.I0(r_4_2_a1_lut6_2_O6[3]),
	.I1(\d_cnst_sn.r_4_0_0 [3]),
	.I2(N_918),
	.I3(N_527_i),
	.I4(N_13),
	.I5(t_1[4]),
	.LO(t_6[4])
);
defparam \d_cnst_sn.reg2_16_11_RNO[4] .INIT=64'hF0004400F0FF44FF;
// @7:103
  LUT6_L \d_cnst_sn.r_4_2_a1_lut6_2_RNI2T8R3[3]  (
	.I0(r_4_2_a1_lut6_2_O6[3]),
	.I1(\d_cnst_sn.r_4_0_0 [3]),
	.I2(N_918),
	.I3(N_527_i),
	.I4(N_13),
	.I5(t_1[4]),
	.LO(r_4_2_a1_lut6_2_RNI2T8R3[3])
);
defparam \d_cnst_sn.r_4_2_a1_lut6_2_RNI2T8R3[3] .INIT=64'h0FFFBBFF0F00BB00;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[8]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_8),
	.I5(un11_reg0_s_8),
	.O(N_1043)
);
defparam \d_cnst_sn.reg0_28_6[8] .INIT=64'hFFFFFF3500CA0000;
// @7:118
  LUT6 un11_r_df20_cZ (
	.I0(N_967),
	.I1(N_935),
	.I2(m_2[20]),
	.I3(m_2[21]),
	.I4(N_13),
	.I5(r_4[21]),
	.O(un11_r_df20)
);
defparam un11_r_df20_cZ.INIT=64'hC300A50000C300A5;
// @7:118
  LUT6 un11_r_lt20_cZ (
	.I0(N_967),
	.I1(N_935),
	.I2(m_2[20]),
	.I3(m_2[21]),
	.I4(N_13),
	.I5(r_4[21]),
	.O(un11_r_lt20)
);
defparam un11_r_lt20_cZ.INIT=64'h30005000FF30FF50;
// @7:151
  LUT6 un26_r_df20_cZ (
	.I0(N_967),
	.I1(N_935),
	.I2(m_2[20]),
	.I3(m_2[21]),
	.I4(N_13),
	.I5(r_4[21]),
	.O(un26_r_df20)
);
defparam un26_r_df20_cZ.INIT=64'hC300A50000C300A5;
// @7:151
  LUT6 un26_r_lt20_cZ (
	.I0(N_967),
	.I1(N_935),
	.I2(m_2[20]),
	.I3(m_2[21]),
	.I4(N_13),
	.I5(r_4[21]),
	.O(un26_r_lt20)
);
defparam un26_r_lt20_cZ.INIT=64'h30005000FF30FF50;
// @7:143
  LUT6 b18_df20_cZ (
	.I0(N_967),
	.I1(N_935),
	.I2(m_2[20]),
	.I3(m_2[21]),
	.I4(N_13),
	.I5(r_4[21]),
	.O(b18_df20)
);
defparam b18_df20_cZ.INIT=64'hC300A50000C300A5;
// @7:143
  LUT6 b18_lt20_cZ (
	.I0(N_967),
	.I1(N_935),
	.I2(m_2[20]),
	.I3(m_2[21]),
	.I4(N_13),
	.I5(r_4[21]),
	.O(b18_lt20)
);
defparam b18_lt20_cZ.INIT=64'h0CFF0AFF000C000A;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[12]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_12),
	.I3(un11_reg0_s_12),
	.O(N_1379)
);
defparam \d_cnst_sn.reg2_16_3[12] .INIT=16'hFD20;
// @7:74
  LUT6_L \d_cnst_sn.reg1_16[0]  (
	.I0(N_513_i),
	.I1(m_2[0]),
	.I2(N_527_i),
	.I3(N_3916),
	.I4(N_1035),
	.I5(t_1[0]),
	.LO(reg1_16[0])
);
defparam \d_cnst_sn.reg1_16[0] .INIT=64'h0044FF44004EFF4E;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28[0]  (
	.I0(N_513_i),
	.I1(m_2[0]),
	.I2(N_527_i),
	.I3(N_3916),
	.I4(N_1035),
	.I5(t_1[0]),
	.LO(reg0_28[0])
);
defparam \d_cnst_sn.reg0_28[0] .INIT=64'h0044FF44004EFF4E;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[15]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_15),
	.I3(un11_reg0_s_15),
	.O(N_1574)
);
defparam \d_cnst_sn.reg2_16_9[15] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[7]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_7),
	.I5(un11_reg0_s_7),
	.O(N_1042)
);
defparam \d_cnst_sn.reg0_28_6[7] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[11]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_11),
	.I5(un11_reg0_s_11),
	.O(N_1046)
);
defparam \d_cnst_sn.reg0_28_6[11] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[13]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_13),
	.I3(un11_reg0_s_13),
	.O(N_1380)
);
defparam \d_cnst_sn.reg2_16_3[13] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[13]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_13),
	.I5(un11_reg0_s_13),
	.O(N_1048)
);
defparam \d_cnst_sn.reg0_28_6[13] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[11]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_11),
	.I3(un11_reg0_s_11),
	.O(N_1378)
);
defparam \d_cnst_sn.reg2_16_3[11] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[10]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_10),
	.I3(un11_reg0_s_10),
	.O(N_1377)
);
defparam \d_cnst_sn.reg2_16_3[10] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[9]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_9),
	.I3(un11_reg0_s_9),
	.O(N_1376)
);
defparam \d_cnst_sn.reg2_16_3[9] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[6]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_6),
	.I3(un11_reg0_s_6),
	.O(N_1373)
);
defparam \d_cnst_sn.reg2_16_3[6] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[3]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_3),
	.I3(un11_reg0_s_3),
	.O(N_1370)
);
defparam \d_cnst_sn.reg2_16_3[3] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[1]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un11_reg0_s_1),
	.I3(un32_reg0_s_1),
	.O(N_1368)
);
defparam \d_cnst_sn.reg2_16_3[1] .INIT=16'hF2D0;
// @7:118
  LUT6 un11_r_df28_cZ (
	.I0(N_943),
	.I1(N_975),
	.I2(m_2[29]),
	.I3(m_2[28]),
	.I4(N_13),
	.I5(r_4[29]),
	.O(un11_r_df28)
);
defparam un11_r_df28_cZ.INIT=64'hA050C0300A050C03;
// @7:118
  LUT6 un11_r_lt28_cZ (
	.I0(N_943),
	.I1(N_975),
	.I2(m_2[29]),
	.I3(m_2[28]),
	.I4(N_13),
	.I5(r_4[29]),
	.O(un11_r_lt28)
);
defparam un11_r_lt28_cZ.INIT=64'h50003000F5F0F3F0;
// @7:151
  LUT6 un26_r_df28_cZ (
	.I0(N_943),
	.I1(N_975),
	.I2(m_2[29]),
	.I3(m_2[28]),
	.I4(N_13),
	.I5(r_4[29]),
	.O(un26_r_df28)
);
defparam un26_r_df28_cZ.INIT=64'hA050C0300A050C03;
// @7:151
  LUT6 un26_r_lt28_cZ (
	.I0(N_943),
	.I1(N_975),
	.I2(m_2[29]),
	.I3(m_2[28]),
	.I4(N_13),
	.I5(r_4[29]),
	.O(un26_r_lt28)
);
defparam un26_r_lt28_cZ.INIT=64'h50003000F5F0F3F0;
// @7:143
  LUT6 b18_df28_cZ (
	.I0(N_943),
	.I1(N_975),
	.I2(m_2[29]),
	.I3(m_2[28]),
	.I4(N_13),
	.I5(r_4[29]),
	.O(b18_df28)
);
defparam b18_df28_cZ.INIT=64'hA050C0300A050C03;
// @7:143
  LUT6 b18_lt28_cZ (
	.I0(N_943),
	.I1(N_975),
	.I2(m_2[29]),
	.I3(m_2[28]),
	.I4(N_13),
	.I5(r_4[29]),
	.O(b18_lt28)
);
defparam b18_lt28_cZ.INIT=64'h0FAF0FCF000A000C;
// @7:118
  LUT6 un11_r_df26_cZ (
	.I0(N_941),
	.I1(N_973),
	.I2(m_2[26]),
	.I3(m_2[27]),
	.I4(N_13),
	.I5(r_4[27]),
	.O(un11_r_df26)
);
defparam un11_r_df26_cZ.INIT=64'hA500C30000A500C3;
// @7:118
  LUT6 un11_r_lt26_cZ (
	.I0(N_941),
	.I1(N_973),
	.I2(m_2[26]),
	.I3(m_2[27]),
	.I4(N_13),
	.I5(r_4[27]),
	.O(un11_r_lt26)
);
defparam un11_r_lt26_cZ.INIT=64'h50003000FF50FF30;
// @7:143
  LUT6 b18_df26_cZ (
	.I0(N_941),
	.I1(N_973),
	.I2(m_2[26]),
	.I3(m_2[27]),
	.I4(N_13),
	.I5(r_4[27]),
	.O(b18_df26)
);
defparam b18_df26_cZ.INIT=64'hA500C30000A500C3;
// @7:151
  LUT6 un26_r_df26_cZ (
	.I0(N_941),
	.I1(N_973),
	.I2(m_2[26]),
	.I3(m_2[27]),
	.I4(N_13),
	.I5(r_4[27]),
	.O(un26_r_df26)
);
defparam un26_r_df26_cZ.INIT=64'hA500C30000A500C3;
// @7:151
  LUT6 un26_r_lt26_cZ (
	.I0(N_941),
	.I1(N_973),
	.I2(m_2[26]),
	.I3(m_2[27]),
	.I4(N_13),
	.I5(r_4[27]),
	.O(un26_r_lt26)
);
defparam un26_r_lt26_cZ.INIT=64'h50003000FF50FF30;
// @7:143
  LUT6 b18_lt26_cZ (
	.I0(N_941),
	.I1(N_973),
	.I2(m_2[26]),
	.I3(m_2[27]),
	.I4(N_13),
	.I5(r_4[27]),
	.O(b18_lt26)
);
defparam b18_lt26_cZ.INIT=64'h0AFF0CFF000A000C;
// @7:118
  LUT6 un11_r_lt24_cZ (
	.I0(N_940),
	.I1(N_972),
	.I2(m_2[24]),
	.I3(m_2[25]),
	.I4(N_13),
	.I5(r_4[24]),
	.O(un11_r_lt24)
);
defparam un11_r_lt24_cZ.INIT=64'h55003300F550F330;
// @7:118
  LUT6 un11_r_df24_cZ (
	.I0(N_940),
	.I1(N_972),
	.I2(m_2[24]),
	.I3(m_2[25]),
	.I4(N_13),
	.I5(r_4[24]),
	.O(un11_r_df24)
);
defparam un11_r_df24_cZ.INIT=64'hA050C0300A050C03;
// @7:143
  LUT6 b18_df24_cZ (
	.I0(N_940),
	.I1(N_972),
	.I2(m_2[24]),
	.I3(m_2[25]),
	.I4(N_13),
	.I5(r_4[24]),
	.O(b18_df24)
);
defparam b18_df24_cZ.INIT=64'hA050C0300A050C03;
// @7:143
  LUT6 b18_lt24_cZ (
	.I0(N_940),
	.I1(N_972),
	.I2(m_2[24]),
	.I3(m_2[25]),
	.I4(N_13),
	.I5(r_4[24]),
	.O(b18_lt24)
);
defparam b18_lt24_cZ.INIT=64'h0AAF0CCF00AA00CC;
// @7:151
  LUT6 un26_r_df24_cZ (
	.I0(N_940),
	.I1(N_972),
	.I2(m_2[24]),
	.I3(m_2[25]),
	.I4(N_13),
	.I5(r_4[24]),
	.O(un26_r_df24)
);
defparam un26_r_df24_cZ.INIT=64'hA050C0300A050C03;
// @7:151
  LUT6 un26_r_lt24_cZ (
	.I0(N_940),
	.I1(N_972),
	.I2(m_2[24]),
	.I3(m_2[25]),
	.I4(N_13),
	.I5(r_4[24]),
	.O(un26_r_lt24)
);
defparam un26_r_lt24_cZ.INIT=64'h55003300F550F330;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11mux_RNO_1[1]  (
	.I0(r_4_2_a0[0]),
	.I1(\d_cnst_sn.r_4_0_0 [0]),
	.I2(N_915),
	.I3(N_527_i),
	.I4(N_13),
	.I5(t_1[1]),
	.LO(t_6[1])
);
defparam \d_cnst_sn.reg2_16_11mux_RNO_1[1] .INIT=64'hF0004400F0FF44FF;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[9]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_9),
	.I5(un11_reg0_s_9),
	.O(N_1044)
);
defparam \d_cnst_sn.reg0_28_6[9] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[1]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un11_reg0_s_1),
	.I5(un32_reg0_s_1),
	.O(N_1036)
);
defparam \d_cnst_sn.reg0_28_6[1] .INIT=64'hFFFF00CAFF350000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[2]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un11_reg0_s_2),
	.I5(un32_reg0_s_2),
	.O(N_1037)
);
defparam \d_cnst_sn.reg0_28_6[2] .INIT=64'hFFFF00CAFF350000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[6]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_6),
	.I5(un11_reg0_s_6),
	.O(N_1041)
);
defparam \d_cnst_sn.reg0_28_6[6] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a4[22]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_22),
	.I5(un11_reg0_s_22),
	.O(reg2_16_11_a4[22])
);
defparam \d_cnst_sn.reg2_16_11_a4[22] .INIT=64'h0000002000100030;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a4[21]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_21),
	.I5(un11_reg0_s_21),
	.O(reg2_16_11_a4[21])
);
defparam \d_cnst_sn.reg2_16_11_a4[21] .INIT=64'h0000002000100030;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a2[17]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_17),
	.I5(un11_reg0_s_17),
	.O(reg2_16_11_a2[17])
);
defparam \d_cnst_sn.reg2_16_11_a2[17] .INIT=64'h000000080004000C;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_1_cZ[20]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.I5(un32_reg0_s_20),
	.O(\d_cnst_sn.reg2_16_1 [20])
);
defparam \d_cnst_sn.reg2_16_1_cZ[20] .INIT=64'hFFFFFFFFFFFFF53F;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[14]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_14),
	.I3(un11_reg0_s_14),
	.O(N_1573)
);
defparam \d_cnst_sn.reg2_16_9[14] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[13]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_13),
	.I3(un11_reg0_s_13),
	.O(N_1572)
);
defparam \d_cnst_sn.reg2_16_9[13] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[12]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_12),
	.I3(un11_reg0_s_12),
	.O(N_1571)
);
defparam \d_cnst_sn.reg2_16_9[12] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[11]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_11),
	.I3(un11_reg0_s_11),
	.O(N_1570)
);
defparam \d_cnst_sn.reg2_16_9[11] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[10]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_10),
	.I3(un11_reg0_s_10),
	.O(N_1569)
);
defparam \d_cnst_sn.reg2_16_9[10] .INIT=16'hFD20;
// @7:47
  LUT5 \d_cnst_sn.addr_20_iv_14_443_i_2_cZ  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_inf_abs0_10[7]),
	.I4(un1_inf_abs0_11[7]),
	.O(\d_cnst_sn.addr_20_iv_14_443_i_2 )
);
defparam \d_cnst_sn.addr_20_iv_14_443_i_2_cZ .INIT=32'h008022A2;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[15]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_15),
	.I3(un11_reg0_s_15),
	.O(N_1382)
);
defparam \d_cnst_sn.reg2_16_3[15] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a4[25]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_25),
	.I5(un11_reg0_s_25),
	.O(reg2_16_11_a4[25])
);
defparam \d_cnst_sn.reg2_16_11_a4[25] .INIT=64'h0000002000100030;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[5]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_5),
	.I3(un11_reg0_s_5),
	.O(N_1372)
);
defparam \d_cnst_sn.reg2_16_3[5] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[16]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_16),
	.I5(un11_reg0_s_16),
	.O(N_1051)
);
defparam \d_cnst_sn.reg0_28_6[16] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[4]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_4),
	.I3(un11_reg0_s_4),
	.O(N_1371)
);
defparam \d_cnst_sn.reg2_16_3[4] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[15]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_15),
	.I5(un11_reg0_s_15),
	.O(N_1050)
);
defparam \d_cnst_sn.reg0_28_6[15] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[17]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_17),
	.I5(un11_reg0_s_17),
	.O(N_1052)
);
defparam \d_cnst_sn.reg0_28_6[17] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[16]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_16),
	.I3(un11_reg0_s_16),
	.O(N_1383)
);
defparam \d_cnst_sn.reg2_16_3[16] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a3[29]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_29),
	.I5(un11_reg0_s_29),
	.O(reg2_16_11_a3[29])
);
defparam \d_cnst_sn.reg2_16_11_a3[29] .INIT=64'h0030001000200000;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a4[24]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_24),
	.I5(un11_reg0_s_24),
	.O(reg2_16_11_a4[24])
);
defparam \d_cnst_sn.reg2_16_11_a4[24] .INIT=64'h0000002000100030;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a2[18]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_18),
	.I5(un11_reg0_s_18),
	.O(reg2_16_11_a2[18])
);
defparam \d_cnst_sn.reg2_16_11_a2[18] .INIT=64'h000000080004000C;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[5]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_5),
	.I3(un11_reg0_s_5),
	.O(N_1564)
);
defparam \d_cnst_sn.reg2_16_9[5] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[10]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_10),
	.I5(un11_reg0_s_10),
	.O(N_1045)
);
defparam \d_cnst_sn.reg0_28_6[10] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[14]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_14),
	.I5(un11_reg0_s_14),
	.O(N_1049)
);
defparam \d_cnst_sn.reg0_28_6[14] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[9]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_9),
	.I3(un11_reg0_s_9),
	.O(N_1568)
);
defparam \d_cnst_sn.reg2_16_9[9] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a2[19]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_19),
	.I5(un11_reg0_s_19),
	.O(reg2_16_11_a2[19])
);
defparam \d_cnst_sn.reg2_16_11_a2[19] .INIT=64'h000000080004000C;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[4]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_4),
	.I5(un11_reg0_s_4),
	.O(N_1039)
);
defparam \d_cnst_sn.reg0_28_6[4] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[18]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_18),
	.I5(un11_reg0_s_18),
	.O(N_1053)
);
defparam \d_cnst_sn.reg0_28_6[18] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[6]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_6),
	.I3(un11_reg0_s_6),
	.O(N_1565)
);
defparam \d_cnst_sn.reg2_16_9[6] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_3[7]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_7),
	.I3(un11_reg0_s_7),
	.O(N_1374)
);
defparam \d_cnst_sn.reg2_16_3[7] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[8]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_8),
	.I3(un11_reg0_s_8),
	.O(N_1567)
);
defparam \d_cnst_sn.reg2_16_9[8] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a4[23]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_23),
	.I5(un11_reg0_s_23),
	.O(reg2_16_11_a4[23])
);
defparam \d_cnst_sn.reg2_16_11_a4[23] .INIT=64'h0000002000100030;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[5]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_5),
	.I5(un11_reg0_s_5),
	.O(N_1040)
);
defparam \d_cnst_sn.reg0_28_6[5] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[3]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_3),
	.I5(un11_reg0_s_3),
	.O(N_1038)
);
defparam \d_cnst_sn.reg0_28_6[3] .INIT=64'hFFFFFF3500CA0000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_6[12]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.I4(un32_reg0_s_12),
	.I5(un11_reg0_s_12),
	.O(N_1047)
);
defparam \d_cnst_sn.reg0_28_6[12] .INIT=64'hFFFFFF3500CA0000;
// @7:47
  LUT4 \d_cnst_sn.reg0_28_11_2228_a6_1_1_cZ  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(reg3_1_1[27]),
	.O(\d_cnst_sn.reg0_28_11_2228_a6_1_1 )
);
defparam \d_cnst_sn.reg0_28_11_2228_a6_1_1_cZ .INIT=16'h0100;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[2]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un11_reg0_s_2),
	.I3(un32_reg0_s_2),
	.O(N_1561)
);
defparam \d_cnst_sn.reg2_16_9[2] .INIT=16'hF2D0;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[25]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_25),
	.I3(un11_reg0_s_25),
	.O(N_1584)
);
defparam \d_cnst_sn.reg2_16_9[25] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[4]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_4),
	.I3(un11_reg0_s_4),
	.O(N_1563)
);
defparam \d_cnst_sn.reg2_16_9[4] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[7]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_7),
	.I3(un11_reg0_s_7),
	.O(N_1566)
);
defparam \d_cnst_sn.reg2_16_9[7] .INIT=16'hFD20;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[3]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un32_reg0_s_3),
	.I3(un11_reg0_s_3),
	.O(N_1562)
);
defparam \d_cnst_sn.reg2_16_9[3] .INIT=16'hFD20;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_2_d[20]  (
	.I0(datai[20]),
	.I1(un3_reg3_s_17),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(inf_abs0_2[27]),
	.I5(inf_abs0_2[28]),
	.O(reg2_16_2_d[20])
);
defparam \d_cnst_sn.reg2_16_2_d[20] .INIT=64'hCCACCCACCCACCC0C;
// @7:74
  LUT4 \d_cnst_sn.reg2_16_9[1]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.I2(un11_reg0_s_1),
	.I3(un32_reg0_s_1),
	.O(N_1560)
);
defparam \d_cnst_sn.reg2_16_9[1] .INIT=16'hF2D0;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[7]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_921),
	.I4(N_953),
	.I5(t_1[7]),
	.LO(t_6[7])
);
defparam \d_cnst_sn.reg2_16_11_RNO[7] .INIT=64'h44400400FFFBBFBB;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[6]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_920),
	.I4(N_952),
	.I5(t_1[6]),
	.LO(t_6[6])
);
defparam \d_cnst_sn.reg2_16_11_RNO[6] .INIT=64'h44400400FFFBBFBB;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[13]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_927),
	.I4(N_959),
	.I5(t_1[13]),
	.LO(t_6[13])
);
defparam \d_cnst_sn.reg2_16_11_RNO[13] .INIT=64'h44400400FFFBBFBB;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[15]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_929),
	.I4(N_961),
	.I5(t_1[15]),
	.LO(t_6[15])
);
defparam \d_cnst_sn.reg2_16_11_RNO[15] .INIT=64'h44400400FFFBBFBB;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[16]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_930),
	.I4(N_962),
	.I5(t_1[16]),
	.LO(t_6[16])
);
defparam \d_cnst_sn.reg2_16_11_RNO[16] .INIT=64'h44400400FFFBBFBB;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[14]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_928),
	.I4(N_960),
	.I5(t_1[14]),
	.LO(t_6[14])
);
defparam \d_cnst_sn.reg2_16_11_RNO[14] .INIT=64'h44400400FFFBBFBB;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_4_a2_0_cZ[20]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_934),
	.I4(N_2722),
	.O(\d_cnst_sn.reg3_17_4_a2_0 [20])
);
defparam \d_cnst_sn.reg3_17_4_a2_0_cZ[20] .INIT=32'h44400400;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[0]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_527_i),
	.I3(N_1335),
	.I4(N_1035),
	.I5(t_1[0]),
	.LO(reg2_16[0])
);
defparam \d_cnst_sn.reg2_16_11[0] .INIT=64'h1100776619087F6E;
// @7:103
  LUT6_L \d_cnst_sn.r_4_1_RNIIQ731[8]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_923),
	.I4(N_955),
	.I5(t_1[9]),
	.LO(r_4_1_RNIIQ731[8])
);
defparam \d_cnst_sn.r_4_1_RNIIQ731[8] .INIT=64'hBBBFFBFF00044044;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[11]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_925),
	.I4(N_957),
	.I5(t_1[11]),
	.LO(t_6[11])
);
defparam \d_cnst_sn.reg2_16_11_RNO[11] .INIT=64'h44400400FFFBBFBB;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[12]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_926),
	.I4(N_958),
	.I5(t_1[12]),
	.LO(t_6[12])
);
defparam \d_cnst_sn.reg2_16_11_RNO[12] .INIT=64'h44400400FFFBBFBB;
// @7:103
  LUT6_L \d_cnst_sn.r_4_1_RNI9K731[5]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_920),
	.I4(N_952),
	.I5(t_1[6]),
	.LO(r_4_1_RNI9K731[5])
);
defparam \d_cnst_sn.r_4_1_RNI9K731[5] .INIT=64'hBBBFFBFF00044044;
// @7:103
  LUT6_L \d_cnst_sn.r_4_1_RNICM731[6]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_921),
	.I4(N_953),
	.I5(t_1[7]),
	.LO(r_4_1_RNICM731[6])
);
defparam \d_cnst_sn.r_4_1_RNICM731[6] .INIT=64'hBBBFFBFF00044044;
// @7:103
  LUT6_L \d_cnst_sn.r_4_1_RNIDBOH1[10]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_925),
	.I4(N_957),
	.I5(t_1[11]),
	.LO(r_4_1_RNIDBOH1[10])
);
defparam \d_cnst_sn.r_4_1_RNIDBOH1[10] .INIT=64'hBBBFFBFF00044044;
// @7:103
  LUT6_L \d_cnst_sn.r_4_1_RNIS3K91[9]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_924),
	.I4(N_956),
	.I5(t_1[10]),
	.LO(r_4_1_RNIS3K91[9])
);
defparam \d_cnst_sn.r_4_1_RNIS3K91[9] .INIT=64'hBBBFFBFF00044044;
// @7:103
  LUT6_L \d_cnst_sn.r_4_1_RNIFO731[7]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_922),
	.I4(N_954),
	.I5(t_1[8]),
	.LO(r_4_1_RNIFO731[7])
);
defparam \d_cnst_sn.r_4_1_RNIFO731[7] .INIT=64'hBBBFFBFF00044044;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_7_a1[17]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[29]),
	.I4(N_931),
	.I5(N_963),
	.O(reg0_28_7_a1[17])
);
defparam \d_cnst_sn.reg0_28_7_a1[17] .INIT=64'h0000002020002020;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[8]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_922),
	.I4(N_954),
	.I5(t_1[8]),
	.LO(t_6[8])
);
defparam \d_cnst_sn.reg2_16_11_RNO[8] .INIT=64'h44400400FFFBBFBB;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[9]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_923),
	.I4(N_955),
	.I5(t_1[9]),
	.LO(t_6[9])
);
defparam \d_cnst_sn.reg2_16_11_RNO[9] .INIT=64'h44400400FFFBBFBB;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_7_a1[18]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(inf_abs0_2[29]),
	.I4(N_932),
	.I5(N_964),
	.O(reg0_28_7_a1[18])
);
defparam \d_cnst_sn.reg0_28_7_a1[18] .INIT=64'h0000002020002020;
// @7:86
  LUT6_L \d_cnst_sn.reg2_16_11_RNO[10]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.I2(inf_abs0_2[29]),
	.I3(N_924),
	.I4(N_956),
	.I5(t_1[10]),
	.LO(t_6[10])
);
defparam \d_cnst_sn.reg2_16_11_RNO[10] .INIT=64'h44400400FFFBBFBB;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_2[23]  (
	.I0(N_7_i),
	.I1(un36_df),
	.I2(un1_b59),
	.I3(un87_df),
	.I4(un32_reg0_s_23),
	.I5(un11_reg0_s_23),
	.LO(N_1742)
);
defparam \d_cnst_sn.reg3_17_2[23] .INIT=64'hFFFFEFFF10000000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_2[24]  (
	.I0(N_7_i),
	.I1(un36_df),
	.I2(un1_b59),
	.I3(un87_df),
	.I4(un32_reg0_s_24),
	.I5(un11_reg0_s_24),
	.LO(N_1743)
);
defparam \d_cnst_sn.reg3_17_2[24] .INIT=64'hFFFFEFFF10000000;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_0[18]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[17]),
	.I4(reg3_1_1[18]),
	.I5(t_1[18]),
	.LO(N_1085)
);
defparam \d_cnst_sn.reg0_28_0[18] .INIT=64'hFDDD2000FFDF2202;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_2[13]  (
	.I0(N_7_i),
	.I1(un36_df),
	.I2(un1_b59),
	.I3(un87_df),
	.I4(un32_reg0_s_13),
	.I5(un11_reg0_s_13),
	.O(N_1732)
);
defparam \d_cnst_sn.reg3_17_2[13] .INIT=64'hFFFFEFFF10000000;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_0[17]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[16]),
	.I4(reg3_1_1[17]),
	.I5(t_1[17]),
	.LO(N_1084)
);
defparam \d_cnst_sn.reg0_28_0[17] .INIT=64'hFDDD2000FFDF2202;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[0]  (
	.I0(datai[0]),
	.I1(m_2[0]),
	.I2(N_1035),
	.I3(un1_cf),
	.I4(N_1810),
	.O(N_1812)
);
defparam \d_cnst_sn.reg3_17_5[0] .INIT=32'hCCAA0F0F;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_2[22]  (
	.I0(N_7_i),
	.I1(un36_df),
	.I2(un1_b59),
	.I3(un87_df),
	.I4(un32_reg0_s_22),
	.I5(un11_reg0_s_22),
	.LO(N_1741)
);
defparam \d_cnst_sn.reg3_17_2[22] .INIT=64'hFFFFEFFF10000000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_2[21]  (
	.I0(N_7_i),
	.I1(un36_df),
	.I2(un1_b59),
	.I3(un87_df),
	.I4(un32_reg0_s_21),
	.I5(un11_reg0_s_21),
	.LO(N_1740)
);
defparam \d_cnst_sn.reg3_17_2[21] .INIT=64'hFFFFEFFF10000000;
// @7:97
  MUXCY_L un3_t_cry_0_cy_cZ (
	.DI(GND),
	.CI(VCC),
	.S(r_4_3_ci[31]),
	.LO(un3_t_cry_0_cy)
);
// @7:97
  LUT6 \d_cnst_sn.r_4_3_ci[31]  (
	.I0(reg0[31]),
	.I1(reg1[31]),
	.I2(reg2[31]),
	.I3(inf_abs0_2[31]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.O(r_4_3_ci[31])
);
defparam \d_cnst_sn.r_4_3_ci[31] .INIT=64'hAA00AAF0AACCAAAA;
// @7:466
  MUXCY_L t_1_cry_0_cy_cZ (
	.DI(GND),
	.CI(VCC),
	.S(r_4_i[31]),
	.LO(t_1_cry_0_cy)
);
  LUT5 \d_cnst_sn.m27  (
	.I0(reg0[2]),
	.I1(reg2[2]),
	.I2(inf_abs0_2[31]),
	.I3(\d_cnst_sn.m19_0_1 ),
	.I4(\d_cnst_sn.m26_0_1 ),
	.O(N_28)
);
defparam \d_cnst_sn.m27 .INIT=32'hACA0AFAA;
// @7:466
  LUT5 un3_t_axb_2_cZ (
	.I0(reg0[2]),
	.I1(reg2[2]),
	.I2(inf_abs0_2[31]),
	.I3(\d_cnst_sn.m19_0_1 ),
	.I4(\d_cnst_sn.m26_0_1 ),
	.O(un3_t_axb_2)
);
defparam un3_t_axb_2_cZ.INIT=32'h535F5055;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_14  (
	.I0(inf_abs0_2[31]),
	.I1(\d_cnst_sn.reg0_28_14_2135_1_a0_2 ),
	.I2(reg3_1_1[30]),
	.I3(\d_cnst_sn.reg0_28_14_0 ),
	.I4(t_1[30]),
	.LO(N_3550)
);
defparam \d_cnst_sn.reg0_28_14 .INIT=32'hFFA0FFEC;
// @7:103
  LUT4 \d_cnst_sn.reg3_17_6_tz[21]  (
	.I0(m_2[21]),
	.I1(\d_cnst_sn.reg3_17_a2_2_0 [21]),
	.I2(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I3(reg3_14_sqmuxa),
	.O(\d_cnst_sn.reg3_17_0_tz [21])
);
defparam \d_cnst_sn.reg3_17_6_tz[21] .INIT=16'hC00A;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28_6_RNIBQPU4[17]  (
	.I0(N_3916),
	.I1(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I2(\d_cnst_sn.reg0_0 [17]),
	.I3(t_1[17]),
	.I4(N_1052),
	.LO(reg0_28[17])
);
defparam \d_cnst_sn.reg0_28_6_RNIBQPU4[17] .INIT=32'hB0F01050;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28_6_RNIGTPU4[18]  (
	.I0(N_3916),
	.I1(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I2(\d_cnst_sn.reg1_0 [18]),
	.I3(t_1[18]),
	.I4(N_1053),
	.LO(reg1_16[18])
);
defparam \d_cnst_sn.reg0_28_6_RNIGTPU4[18] .INIT=32'hB0F01050;
// @7:74
  LUT1_L \state_RNO[0]  (
	.I0(state[0]),
	.LO(state_i[0])
);
defparam \state_RNO[0] .INIT=2'h1;
// @7:74
  LUT2 un1_inf_abs0_0_s_19_RNO (
	.I0(reg1[19]),
	.I1(inf_abs0_2[19]),
	.O(un1_inf_abs0_0_axb_19)
);
defparam un1_inf_abs0_0_s_19_RNO.INIT=4'h6;
// @7:74
  LUT2 un1_inf_abs0_s_19_RNO (
	.I0(reg2[19]),
	.I1(inf_abs0_2[19]),
	.O(un1_inf_abs0_axb_19)
);
defparam un1_inf_abs0_s_19_RNO.INIT=4'h6;
  LUT2 \d_cnst_sn.m2  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[30]),
	.O(N_3_0)
);
defparam \d_cnst_sn.m2 .INIT=4'h4;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[8]  (
	.I0(datai[8]),
	.I1(state[0]),
	.I2(inf_abs0_2[8]),
	.LO(ir_3[8])
);
defparam \d_cnst_sn.ir_3[8] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[16]  (
	.I0(datai[16]),
	.I1(state[0]),
	.I2(inf_abs0_2[16]),
	.LO(ir_3[16])
);
defparam \d_cnst_sn.ir_3[16] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[3]  (
	.I0(datai[3]),
	.I1(state[0]),
	.I2(inf_abs0_2[3]),
	.LO(ir_3[3])
);
defparam \d_cnst_sn.ir_3[3] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[0]  (
	.I0(datai[0]),
	.I1(state[0]),
	.I2(inf_abs0_2[0]),
	.LO(ir_3[0])
);
defparam \d_cnst_sn.ir_3[0] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[27]  (
	.I0(datai[27]),
	.I1(state[0]),
	.I2(inf_abs0_2[27]),
	.LO(ir_3[27])
);
defparam \d_cnst_sn.ir_3[27] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[23]  (
	.I0(datai[23]),
	.I1(state[0]),
	.I2(inf_abs0_2[23]),
	.LO(ir_3[23])
);
defparam \d_cnst_sn.ir_3[23] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[26]  (
	.I0(datai[26]),
	.I1(state[0]),
	.I2(inf_abs0_2[26]),
	.LO(ir_3[26])
);
defparam \d_cnst_sn.ir_3[26] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[5]  (
	.I0(datai[5]),
	.I1(state[0]),
	.I2(inf_abs0_2[5]),
	.LO(ir_3[5])
);
defparam \d_cnst_sn.ir_3[5] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[2]  (
	.I0(datai[2]),
	.I1(state[0]),
	.I2(inf_abs0_2[2]),
	.LO(ir_3[2])
);
defparam \d_cnst_sn.ir_3[2] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[18]  (
	.I0(datai[18]),
	.I1(state[0]),
	.I2(inf_abs0_2[18]),
	.LO(ir_3[18])
);
defparam \d_cnst_sn.ir_3[18] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[19]  (
	.I0(datai[19]),
	.I1(state[0]),
	.I2(inf_abs0_2[19]),
	.LO(ir_3[19])
);
defparam \d_cnst_sn.ir_3[19] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[10]  (
	.I0(datai[10]),
	.I1(state[0]),
	.I2(inf_abs0_2[10]),
	.LO(ir_3[10])
);
defparam \d_cnst_sn.ir_3[10] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[9]  (
	.I0(datai[9]),
	.I1(state[0]),
	.I2(inf_abs0_2[9]),
	.LO(ir_3[9])
);
defparam \d_cnst_sn.ir_3[9] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[6]  (
	.I0(datai[6]),
	.I1(state[0]),
	.I2(inf_abs0_2[6]),
	.LO(ir_3[6])
);
defparam \d_cnst_sn.ir_3[6] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[4]  (
	.I0(datai[4]),
	.I1(state[0]),
	.I2(inf_abs0_2[4]),
	.LO(ir_3[4])
);
defparam \d_cnst_sn.ir_3[4] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[22]  (
	.I0(datai[22]),
	.I1(state[0]),
	.I2(inf_abs0_2[22]),
	.LO(ir_3[22])
);
defparam \d_cnst_sn.ir_3[22] .INIT=8'hE2;
// @7:47
  LUT3 \d_cnst_sn.r_4_3_21_1130_i_m4  (
	.I0(reg1[19]),
	.I1(un3_reg3_s_16),
	.I2(inf_abs0_2[30]),
	.O(N_2722)
);
defparam \d_cnst_sn.r_4_3_21_1130_i_m4 .INIT=8'hCA;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[21]  (
	.I0(datai[21]),
	.I1(state[0]),
	.I2(inf_abs0_2[21]),
	.LO(ir_3[21])
);
defparam \d_cnst_sn.ir_3[21] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[1]  (
	.I0(datai[1]),
	.I1(state[0]),
	.I2(inf_abs0_2[1]),
	.LO(ir_3[1])
);
defparam \d_cnst_sn.ir_3[1] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[7]  (
	.I0(datai[7]),
	.I1(state[0]),
	.I2(inf_abs0_2[7]),
	.LO(ir_3[7])
);
defparam \d_cnst_sn.ir_3[7] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[25]  (
	.I0(datai[25]),
	.I1(state[0]),
	.I2(inf_abs0_2[25]),
	.LO(ir_3[25])
);
defparam \d_cnst_sn.ir_3[25] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[24]  (
	.I0(datai[24]),
	.I1(state[0]),
	.I2(inf_abs0_2[24]),
	.LO(ir_3[24])
);
defparam \d_cnst_sn.ir_3[24] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[29]  (
	.I0(datai[29]),
	.I1(state[0]),
	.I2(inf_abs0_2[29]),
	.LO(ir_3[29])
);
defparam \d_cnst_sn.ir_3[29] .INIT=8'hE2;
// @7:74
  LUT3_L \d_cnst_sn.ir_3[11]  (
	.I0(datai[11]),
	.I1(state[0]),
	.I2(inf_abs0_2[11]),
	.LO(ir_3[11])
);
defparam \d_cnst_sn.ir_3[11] .INIT=8'hE2;
// @7:97
  LUT3 \d_cnst_sn.r_4_2_a0[0]  (
	.I0(reg3[0]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[30]),
	.O(r_4_2_a0[0])
);
defparam \d_cnst_sn.r_4_2_a0[0] .INIT=8'h10;
// @7:97
  LUT3 \d_cnst_sn.r_4_2_a0[1]  (
	.I0(reg3[1]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[30]),
	.O(r_4_2_a0[1])
);
defparam \d_cnst_sn.r_4_2_a0[1] .INIT=8'h10;
// @7:97
  LUT3 \d_cnst_sn.r_4_0_0_0[0]  (
	.I0(reg1[0]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[30]),
	.O(\d_cnst_sn.r_4_0_0 [0])
);
defparam \d_cnst_sn.r_4_0_0_0[0] .INIT=8'hBA;
// @7:97
  LUT3 \d_cnst_sn.r_4_0_0_cZ[1]  (
	.I0(reg1[1]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[30]),
	.O(\d_cnst_sn.r_4_0_0 [1])
);
defparam \d_cnst_sn.r_4_0_0_cZ[1] .INIT=8'hBA;
// @7:106
  LUT3 \d_cnst_sn.m7_0  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.O(m7)
);
defparam \d_cnst_sn.m7_0 .INIT=8'hAB;
// @7:83
  LUT2 inf_abs0_2_axb_30_cZ (
	.I0(ir[30]),
	.I1(ir[31]),
	.O(inf_abs0_2_axb_30)
);
defparam inf_abs0_2_axb_30_cZ.INIT=4'h6;
// @7:92
  LUT2 \un9_cf_1.SUM0  (
	.I0(inf_abs0_2[23]),
	.I1(inf_abs0_2[31]),
	.O(N_7_i)
);
defparam \un9_cf_1.SUM0 .INIT=4'h2;
  LUT2 \d_cnst_sn.m12  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.O(N_13)
);
defparam \d_cnst_sn.m12 .INIT=4'hB;
// @7:90
  LUT2 \d_cnst_sn.SUM3  (
	.I0(inf_abs0_2[22]),
	.I1(inf_abs0_2[31]),
	.O(N_514_i)
);
defparam \d_cnst_sn.SUM3 .INIT=4'h2;
// @7:90
  LUT2 \d_cnst_sn.SUM2_0  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.O(N_513_i)
);
defparam \d_cnst_sn.SUM2_0 .INIT=4'h2;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[11]  (
	.I0(reg0[11]),
	.I1(reg2[11]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_926)
);
defparam \d_cnst_sn.r_4_1[11] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[26]  (
	.I0(reg0[26]),
	.I1(reg2[26]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_941)
);
defparam \d_cnst_sn.r_4_1[26] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[11]  (
	.I0(reg1[11]),
	.I1(un3_reg3_s_8),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_958)
);
defparam \d_cnst_sn.r_4_2[11] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[26]  (
	.I0(reg1[26]),
	.I1(un3_reg3_s_23),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_973)
);
defparam \d_cnst_sn.r_4_2[26] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[28]  (
	.I0(reg0[28]),
	.I1(reg2[28]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_943)
);
defparam \d_cnst_sn.r_4_1[28] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[28]  (
	.I0(reg1[28]),
	.I1(un3_reg3_s_25),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_975)
);
defparam \d_cnst_sn.r_4_2[28] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[25]  (
	.I0(reg0[25]),
	.I1(reg2[25]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_940)
);
defparam \d_cnst_sn.r_4_1[25] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[25]  (
	.I0(reg1[25]),
	.I1(un3_reg3_s_22),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_972)
);
defparam \d_cnst_sn.r_4_2[25] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[13]  (
	.I0(reg0[13]),
	.I1(reg2[13]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_928)
);
defparam \d_cnst_sn.r_4_1[13] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[13]  (
	.I0(reg1[13]),
	.I1(un3_reg3_s_10),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_960)
);
defparam \d_cnst_sn.r_4_2[13] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[16]  (
	.I0(reg0[16]),
	.I1(reg2[16]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_931)
);
defparam \d_cnst_sn.r_4_1[16] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[16]  (
	.I0(reg1[16]),
	.I1(un3_reg3_s_13),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_963)
);
defparam \d_cnst_sn.r_4_2[16] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[14]  (
	.I0(reg0[14]),
	.I1(reg2[14]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_929)
);
defparam \d_cnst_sn.r_4_1[14] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[14]  (
	.I0(reg1[14]),
	.I1(un3_reg3_s_11),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_961)
);
defparam \d_cnst_sn.r_4_2[14] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[10]  (
	.I0(reg0[10]),
	.I1(reg2[10]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_925)
);
defparam \d_cnst_sn.r_4_1[10] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[10]  (
	.I0(reg1[10]),
	.I1(un3_reg3_s_7),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_957)
);
defparam \d_cnst_sn.r_4_2[10] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[9]  (
	.I0(reg0[9]),
	.I1(reg2[9]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_924)
);
defparam \d_cnst_sn.r_4_1[9] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[9]  (
	.I0(reg1[9]),
	.I1(un3_reg3_s_6),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_956)
);
defparam \d_cnst_sn.r_4_2[9] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[7]  (
	.I0(reg0[7]),
	.I1(reg2[7]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_922)
);
defparam \d_cnst_sn.r_4_1[7] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[8]  (
	.I0(reg0[8]),
	.I1(reg2[8]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_923)
);
defparam \d_cnst_sn.r_4_1[8] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[7]  (
	.I0(reg1[7]),
	.I1(un3_reg3_s_4),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_954)
);
defparam \d_cnst_sn.r_4_2[7] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[8]  (
	.I0(reg1[8]),
	.I1(un3_reg3_s_5),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_955)
);
defparam \d_cnst_sn.r_4_2[8] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[21]  (
	.I0(reg0[21]),
	.I1(reg2[21]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_936)
);
defparam \d_cnst_sn.r_4_1[21] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[21]  (
	.I0(reg1[21]),
	.I1(un3_reg3_s_18),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_968)
);
defparam \d_cnst_sn.r_4_2[21] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[20]  (
	.I0(reg0[20]),
	.I1(reg2[20]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_935)
);
defparam \d_cnst_sn.r_4_1[20] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[20]  (
	.I0(reg1[20]),
	.I1(un3_reg3_s_17),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_967)
);
defparam \d_cnst_sn.r_4_2[20] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[15]  (
	.I0(reg0[15]),
	.I1(reg2[15]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_930)
);
defparam \d_cnst_sn.r_4_1[15] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[17]  (
	.I0(reg0[17]),
	.I1(reg2[17]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_932)
);
defparam \d_cnst_sn.r_4_1[17] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[15]  (
	.I0(reg1[15]),
	.I1(un3_reg3_s_12),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_962)
);
defparam \d_cnst_sn.r_4_2[15] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[17]  (
	.I0(reg1[17]),
	.I1(un3_reg3_s_14),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_964)
);
defparam \d_cnst_sn.r_4_2[17] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[5]  (
	.I0(reg0[5]),
	.I1(reg2[5]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_920)
);
defparam \d_cnst_sn.r_4_1[5] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[5]  (
	.I0(reg1[5]),
	.I1(un3_reg3_s_2),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_952)
);
defparam \d_cnst_sn.r_4_2[5] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[27]  (
	.I0(reg0[27]),
	.I1(reg2[27]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_942)
);
defparam \d_cnst_sn.r_4_1[27] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[27]  (
	.I0(reg1[27]),
	.I1(un3_reg3_s_24),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_974)
);
defparam \d_cnst_sn.r_4_2[27] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[18]  (
	.I0(reg0[18]),
	.I1(reg2[18]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_933)
);
defparam \d_cnst_sn.r_4_1[18] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[18]  (
	.I0(reg1[18]),
	.I1(un3_reg3_s_15),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_965)
);
defparam \d_cnst_sn.r_4_2[18] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[22]  (
	.I0(reg0[22]),
	.I1(reg2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_937)
);
defparam \d_cnst_sn.r_4_1[22] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[22]  (
	.I0(reg1[22]),
	.I1(un3_reg3_s_19),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_969)
);
defparam \d_cnst_sn.r_4_2[22] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[12]  (
	.I0(reg0[12]),
	.I1(reg2[12]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_927)
);
defparam \d_cnst_sn.r_4_1[12] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[12]  (
	.I0(reg1[12]),
	.I1(un3_reg3_s_9),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_959)
);
defparam \d_cnst_sn.r_4_2[12] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[6]  (
	.I0(reg0[6]),
	.I1(reg2[6]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_921)
);
defparam \d_cnst_sn.r_4_1[6] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[6]  (
	.I0(reg1[6]),
	.I1(un3_reg3_s_3),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_953)
);
defparam \d_cnst_sn.r_4_2[6] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[19]  (
	.I0(reg0[19]),
	.I1(reg2[19]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_934)
);
defparam \d_cnst_sn.r_4_1[19] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[23]  (
	.I0(reg1[23]),
	.I1(un3_reg3_s_20),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_970)
);
defparam \d_cnst_sn.r_4_2[23] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[23]  (
	.I0(reg0[23]),
	.I1(reg2[23]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_938)
);
defparam \d_cnst_sn.r_4_1[23] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_2[24]  (
	.I0(reg1[24]),
	.I1(un3_reg3_s_21),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_971)
);
defparam \d_cnst_sn.r_4_2[24] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4_1[24]  (
	.I0(reg0[24]),
	.I1(reg2[24]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_939)
);
defparam \d_cnst_sn.r_4_1[24] .INIT=16'hACAA;
  LUT4 \d_cnst_sn.m19_0_1_cZ  (
	.I0(reg1[2]),
	.I1(reg3[2]),
	.I2(inf_abs0_2[29]),
	.I3(inf_abs0_2[30]),
	.O(\d_cnst_sn.m19_0_1 )
);
defparam \d_cnst_sn.m19_0_1_cZ .INIT=16'hCFA0;
  LUT4 \d_cnst_sn.m26_0_1_cZ  (
	.I0(reg1[2]),
	.I1(reg3[2]),
	.I2(inf_abs0_2[29]),
	.I3(inf_abs0_2[30]),
	.O(\d_cnst_sn.m26_0_1 )
);
defparam \d_cnst_sn.m26_0_1_cZ .INIT=16'h3F50;
// @7:97
  LUT4 \d_cnst_sn.r_4_0_0_0[3]  (
	.I0(reg1[3]),
	.I1(reg3[3]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(\d_cnst_sn.r_4_0_0 [3])
);
defparam \d_cnst_sn.r_4_0_0_0[3] .INIT=16'hA3AF;
// @7:97
  LUT4 \d_cnst_sn.r_4_0_0_0[4]  (
	.I0(reg1[4]),
	.I1(un3_reg3_s_1),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(\d_cnst_sn.r_4_0_0 [4])
);
defparam \d_cnst_sn.r_4_0_0_0[4] .INIT=16'hACAF;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_26  (
	.I0(m_2[22]),
	.I1(m_2[23]),
	.I2(m_2[21]),
	.I3(r_4[21]),
	.I4(r_4[23]),
	.I5(r_4[22]),
	.O(un14_r_0_N_56)
);
defparam \d_cnst_sn.un14_r_0_I_26 .INIT=64'h8008200240041001;
// @7:47
  LUT5 \d_cnst_sn.addr_20_iv_0_1025_i_a6_3  (
	.I0(state[0]),
	.I1(inf_abs0_2[24]),
	.I2(inf_abs0_2[23]),
	.I3(inf_abs0_2[25]),
	.I4(inf_abs0_2[26]),
	.O(N_2641)
);
defparam \d_cnst_sn.addr_20_iv_0_1025_i_a6_3 .INIT=32'h08000000;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_50  (
	.I0(m_2[24]),
	.I1(m_2[25]),
	.I2(m_2[26]),
	.I3(r_4[24]),
	.I4(r_4[25]),
	.I5(r_4[26]),
	.O(un14_r_0_N_35)
);
defparam \d_cnst_sn.un14_r_0_I_50 .INIT=64'h8040201008040201;
// @7:97
  LUT4 \d_cnst_sn.r_4[0]  (
	.I0(reg0[0]),
	.I1(reg2[0]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_915)
);
defparam \d_cnst_sn.r_4[0] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4[1]  (
	.I0(reg0[1]),
	.I1(reg2[1]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_916)
);
defparam \d_cnst_sn.r_4[1] .INIT=16'hACAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_6_1508_i_m2  (
	.I0(reg0[29]),
	.I1(reg1[29]),
	.I2(reg2[29]),
	.I3(un3_reg3_cry_25),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_6_1508_i_m2)
);
defparam \d_cnst_sn.r_4_3_6_1508_i_m2 .INIT=64'hFF00F0F0CCCCAAAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_5_1534_i_m2  (
	.I0(reg1[28]),
	.I1(reg0[28]),
	.I2(reg2[28]),
	.I3(un3_reg3_s_25),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_5_1534_i_m2)
);
defparam \d_cnst_sn.r_4_3_5_1534_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_1_1638_i_m2  (
	.I0(reg0[24]),
	.I1(reg2[24]),
	.I2(reg1[24]),
	.I3(un3_reg3_s_21),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_1_1638_i_m2)
);
defparam \d_cnst_sn.r_4_3_1_1638_i_m2 .INIT=64'hFF00CCCCF0F0AAAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_18_1208_i_m2  (
	.I0(reg1[16]),
	.I1(reg0[16]),
	.I2(reg2[16]),
	.I3(un3_reg3_s_13),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_18_1208_i_m2)
);
defparam \d_cnst_sn.r_4_3_18_1208_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_15_1286_i_m2  (
	.I0(reg1[13]),
	.I1(reg0[13]),
	.I2(reg2[13]),
	.I3(un3_reg3_s_10),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_15_1286_i_m2)
);
defparam \d_cnst_sn.r_4_3_15_1286_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_13_1338_i_m2  (
	.I0(reg1[11]),
	.I1(reg0[11]),
	.I2(reg2[11]),
	.I3(un3_reg3_s_8),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_13_1338_i_m2)
);
defparam \d_cnst_sn.r_4_3_13_1338_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_19_1182_i_m2  (
	.I0(reg1[17]),
	.I1(reg0[17]),
	.I2(reg2[17]),
	.I3(un3_reg3_s_14),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_19_1182_i_m2)
);
defparam \d_cnst_sn.r_4_3_19_1182_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_14_1312_i_m2  (
	.I0(reg1[12]),
	.I1(reg0[12]),
	.I2(reg2[12]),
	.I3(un3_reg3_s_9),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_14_1312_i_m2)
);
defparam \d_cnst_sn.r_4_3_14_1312_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_12_1364_i_m2  (
	.I0(reg1[10]),
	.I1(reg0[10]),
	.I2(reg2[10]),
	.I3(un3_reg3_s_7),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_12_1364_i_m2)
);
defparam \d_cnst_sn.r_4_3_12_1364_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_3_1586_i_m2  (
	.I0(reg1[26]),
	.I1(reg0[26]),
	.I2(reg2[26]),
	.I3(un3_reg3_s_23),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_3_1586_i_m2)
);
defparam \d_cnst_sn.r_4_3_3_1586_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_16_1260_i_m2  (
	.I0(reg1[14]),
	.I1(reg0[14]),
	.I2(reg2[14]),
	.I3(un3_reg3_s_11),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_16_1260_i_m2)
);
defparam \d_cnst_sn.r_4_3_16_1260_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_11_1390_i_m2  (
	.I0(reg1[9]),
	.I1(reg0[9]),
	.I2(reg2[9]),
	.I3(un3_reg3_s_6),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_11_1390_i_m2)
);
defparam \d_cnst_sn.r_4_3_11_1390_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_30_680_i_m2  (
	.I0(reg1[6]),
	.I1(reg0[6]),
	.I2(reg2[6]),
	.I3(un3_reg3_s_3),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_30_680_i_m2)
);
defparam \d_cnst_sn.r_4_3_30_680_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_10_1416_i_m2  (
	.I0(reg1[8]),
	.I1(reg0[8]),
	.I2(reg2[8]),
	.I3(un3_reg3_s_5),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_10_1416_i_m2)
);
defparam \d_cnst_sn.r_4_3_10_1416_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_9_1442_i_m2  (
	.I0(reg1[7]),
	.I1(reg0[7]),
	.I2(reg2[7]),
	.I3(un3_reg3_s_4),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_9_1442_i_m2)
);
defparam \d_cnst_sn.r_4_3_9_1442_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_0_1664_i_m2  (
	.I0(reg0[23]),
	.I1(reg2[23]),
	.I2(reg1[23]),
	.I3(un3_reg3_s_20),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_0_1664_i_m2)
);
defparam \d_cnst_sn.r_4_3_0_1664_i_m2 .INIT=64'hFF00CCCCF0F0AAAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_22_1104_i_m2  (
	.I0(reg0[20]),
	.I1(reg2[20]),
	.I2(reg1[20]),
	.I3(un3_reg3_s_17),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_22_1104_i_m2)
);
defparam \d_cnst_sn.r_4_3_22_1104_i_m2 .INIT=64'hFF00CCCCF0F0AAAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_25_810_i_m2  (
	.I0(reg0[1]),
	.I1(reg2[1]),
	.I2(reg1[1]),
	.I3(reg3[1]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_25_810_i_m2)
);
defparam \d_cnst_sn.r_4_3_25_810_i_m2 .INIT=64'hFF00CCCCF0F0AAAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_17_1234_i_m2  (
	.I0(reg1[15]),
	.I1(reg0[15]),
	.I2(reg2[15]),
	.I3(un3_reg3_s_12),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_17_1234_i_m2)
);
defparam \d_cnst_sn.r_4_3_17_1234_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_29_706_i_m2  (
	.I0(reg1[5]),
	.I1(reg0[5]),
	.I2(reg2[5]),
	.I3(un3_reg3_s_2),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_29_706_i_m2)
);
defparam \d_cnst_sn.r_4_3_29_706_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_24_836_i_m2  (
	.I0(reg0[0]),
	.I1(reg2[0]),
	.I2(reg1[0]),
	.I3(reg3[0]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_24_836_i_m2)
);
defparam \d_cnst_sn.r_4_3_24_836_i_m2 .INIT=64'hFF00CCCCF0F0AAAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_4_1560_i_m2  (
	.I0(reg0[27]),
	.I1(reg2[27]),
	.I2(reg1[27]),
	.I3(un3_reg3_s_24),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_4_1560_i_m2)
);
defparam \d_cnst_sn.r_4_3_4_1560_i_m2 .INIT=64'hFF00CCCCF0F0AAAA;
// @7:105
  LUT4 \d_cnst_sn.m_2[29]  (
	.I0(datai[29]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[29])
);
defparam \d_cnst_sn.m_2[29] .INIT=16'h2220;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_20_1156_i_m2  (
	.I0(reg1[18]),
	.I1(reg0[18]),
	.I2(reg2[18]),
	.I3(un3_reg3_s_15),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_20_1156_i_m2)
);
defparam \d_cnst_sn.r_4_3_20_1156_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_1690_i_m2  (
	.I0(reg0[22]),
	.I1(reg2[22]),
	.I2(reg1[22]),
	.I3(un3_reg3_s_19),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_1690_i_m2)
);
defparam \d_cnst_sn.r_4_3_1690_i_m2 .INIT=64'hFF00CCCCF0F0AAAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_28_732_i_m2  (
	.I0(reg0[4]),
	.I1(reg2[4]),
	.I2(reg1[4]),
	.I3(un3_reg3_s_1),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_28_732_i_m2)
);
defparam \d_cnst_sn.r_4_3_28_732_i_m2 .INIT=64'hFF00CCCCF0F0AAAA;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_2_1612_i_m2  (
	.I0(reg1[25]),
	.I1(reg0[25]),
	.I2(reg2[25]),
	.I3(un3_reg3_s_22),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_2_1612_i_m2)
);
defparam \d_cnst_sn.r_4_3_2_1612_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_23_1078_i_m2  (
	.I0(reg1[21]),
	.I1(reg0[21]),
	.I2(reg2[21]),
	.I3(un3_reg3_s_18),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_23_1078_i_m2)
);
defparam \d_cnst_sn.r_4_3_23_1078_i_m2 .INIT=64'hFF00F0F0AAAACCCC;
// @7:47
  LUT6_L \d_cnst_sn.r_4_3_27_758_i_m2  (
	.I0(reg0[3]),
	.I1(reg2[3]),
	.I2(reg1[3]),
	.I3(reg3[3]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(r_4_3_27_758_i_m2)
);
defparam \d_cnst_sn.r_4_3_27_758_i_m2 .INIT=64'h00FFCCCCF0F0AAAA;
// @7:227
  LUT3 \d_cnst_sn.un1_reg0_0_sqmuxa_1_i_o4  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[31]),
	.O(N_1901)
);
defparam \d_cnst_sn.un1_reg0_0_sqmuxa_1_i_o4 .INIT=8'h0E;
// @7:105
  LUT5 \d_cnst_sn.m_2[5]  (
	.I0(datai[5]),
	.I1(inf_abs0_2[5]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[5])
);
defparam \d_cnst_sn.m_2[5] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[8]  (
	.I0(datai[8]),
	.I1(inf_abs0_2[8]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[8])
);
defparam \d_cnst_sn.m_2[8] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[15]  (
	.I0(datai[15]),
	.I1(inf_abs0_2[15]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[15])
);
defparam \d_cnst_sn.m_2[15] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[16]  (
	.I0(datai[16]),
	.I1(inf_abs0_2[16]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[16])
);
defparam \d_cnst_sn.m_2[16] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[3]  (
	.I0(datai[3]),
	.I1(inf_abs0_2[3]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[3])
);
defparam \d_cnst_sn.m_2[3] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[1]  (
	.I0(datai[1]),
	.I1(inf_abs0_2[1]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[1])
);
defparam \d_cnst_sn.m_2[1] .INIT=32'hCACACACC;
// @7:47
  LUT5_L \d_cnst_sn.r_4_3_8_1467  (
	.I0(reg0[31]),
	.I1(reg1[31]),
	.I2(reg2[31]),
	.I3(inf_abs0_2[29]),
	.I4(inf_abs0_2[30]),
	.LO(r_4_3_8_1467)
);
defparam \d_cnst_sn.r_4_3_8_1467 .INIT=32'h00F0CCAA;
// @7:105
  LUT5 \d_cnst_sn.m_2[13]  (
	.I0(datai[13]),
	.I1(inf_abs0_2[13]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[13])
);
defparam \d_cnst_sn.m_2[13] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[19]  (
	.I0(datai[19]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[19])
);
defparam \d_cnst_sn.m_2[19] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[14]  (
	.I0(datai[14]),
	.I1(inf_abs0_2[14]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[14])
);
defparam \d_cnst_sn.m_2[14] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[18]  (
	.I0(datai[18]),
	.I1(inf_abs0_2[18]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[18])
);
defparam \d_cnst_sn.m_2[18] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[12]  (
	.I0(datai[12]),
	.I1(inf_abs0_2[12]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[12])
);
defparam \d_cnst_sn.m_2[12] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[17]  (
	.I0(datai[17]),
	.I1(inf_abs0_2[17]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[17])
);
defparam \d_cnst_sn.m_2[17] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[10]  (
	.I0(datai[10]),
	.I1(inf_abs0_2[10]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[10])
);
defparam \d_cnst_sn.m_2[10] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[11]  (
	.I0(datai[11]),
	.I1(inf_abs0_2[11]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[11])
);
defparam \d_cnst_sn.m_2[11] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[9]  (
	.I0(datai[9]),
	.I1(inf_abs0_2[9]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[9])
);
defparam \d_cnst_sn.m_2[9] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[2]  (
	.I0(datai[2]),
	.I1(inf_abs0_2[2]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[2])
);
defparam \d_cnst_sn.m_2[2] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[6]  (
	.I0(datai[6]),
	.I1(inf_abs0_2[6]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[6])
);
defparam \d_cnst_sn.m_2[6] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[7]  (
	.I0(datai[7]),
	.I1(inf_abs0_2[7]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[7])
);
defparam \d_cnst_sn.m_2[7] .INIT=32'hCACACACC;
// @7:105
  LUT5 \d_cnst_sn.m_2[4]  (
	.I0(datai[4]),
	.I1(inf_abs0_2[4]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[4])
);
defparam \d_cnst_sn.m_2[4] .INIT=32'hCACACACC;
// @7:47
  LUT5_L \d_cnst_sn.addr_20_iv_18_335_i_1_cZ  (
	.I0(reg3[11]),
	.I1(state[0]),
	.I2(inf_abs0_2[11]),
	.I3(inf_abs0_2[28]),
	.I4(N_2641),
	.LO(\d_cnst_sn.addr_20_iv_18_335_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_18_335_i_1_cZ .INIT=32'hFFFF111D;
// @7:47
  LUT5_L \d_cnst_sn.addr_20_iv_13_470_i_1_cZ  (
	.I0(reg3[6]),
	.I1(state[0]),
	.I2(inf_abs0_2[6]),
	.I3(inf_abs0_2[28]),
	.I4(N_2641),
	.LO(\d_cnst_sn.addr_20_iv_13_470_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_13_470_i_1_cZ .INIT=32'hFFFF111D;
// @7:47
  LUT5_L \d_cnst_sn.addr_20_iv_17_362_i_1_cZ  (
	.I0(reg3[10]),
	.I1(state[0]),
	.I2(inf_abs0_2[10]),
	.I3(inf_abs0_2[28]),
	.I4(N_2641),
	.LO(\d_cnst_sn.addr_20_iv_17_362_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_17_362_i_1_cZ .INIT=32'hFFFF111D;
// @7:47
  LUT5_L \d_cnst_sn.addr_20_iv_15_416_i_1_cZ  (
	.I0(reg3[8]),
	.I1(state[0]),
	.I2(inf_abs0_2[8]),
	.I3(inf_abs0_2[28]),
	.I4(N_2641),
	.LO(\d_cnst_sn.addr_20_iv_15_416_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_15_416_i_1_cZ .INIT=32'hFFFF111D;
// @7:47
  LUT5_L \d_cnst_sn.addr_20_iv_10_562_i_1_cZ  (
	.I0(reg3[3]),
	.I1(state[0]),
	.I2(inf_abs0_2[3]),
	.I3(inf_abs0_2[28]),
	.I4(N_2641),
	.LO(\d_cnst_sn.addr_20_iv_10_562_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_10_562_i_1_cZ .INIT=32'hFFFF111D;
// @7:47
  LUT5_L \d_cnst_sn.addr_20_iv_12_497_i_1_cZ  (
	.I0(reg3[5]),
	.I1(state[0]),
	.I2(inf_abs0_2[5]),
	.I3(inf_abs0_2[28]),
	.I4(N_2641),
	.LO(\d_cnst_sn.addr_20_iv_12_497_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_12_497_i_1_cZ .INIT=32'hFFFF111D;
// @7:47
  LUT5_L \d_cnst_sn.addr_20_iv_16_389_i_1_cZ  (
	.I0(reg3[9]),
	.I1(state[0]),
	.I2(inf_abs0_2[9]),
	.I3(inf_abs0_2[28]),
	.I4(N_2641),
	.LO(\d_cnst_sn.addr_20_iv_16_389_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_16_389_i_1_cZ .INIT=32'hFFFF111D;
// @7:47
  LUT6 \d_cnst_sn.addr_20_iv_8_627_i_1_cZ  (
	.I0(reg3[1]),
	.I1(state[0]),
	.I2(inf_abs0_2[1]),
	.I3(un1_inf_abs0_11[1]),
	.I4(inf_abs0_2[27]),
	.I5(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_8_627_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_8_627_i_1_cZ .INIT=64'h111111DD1D1D1DDD;
// @7:97
  LUT4 \d_cnst_sn.r_4[4]  (
	.I0(reg0[4]),
	.I1(reg2[4]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_919)
);
defparam \d_cnst_sn.r_4[4] .INIT=16'hACAA;
// @7:97
  LUT4 \d_cnst_sn.r_4[3]  (
	.I0(reg0[3]),
	.I1(reg2[3]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[30]),
	.O(N_918)
);
defparam \d_cnst_sn.r_4[3] .INIT=16'hACAA;
// @7:74
  LUT5 \d_cnst_sn.un1_state_1_1_o6_0  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.O(N_1890)
);
defparam \d_cnst_sn.un1_state_1_1_o6_0 .INIT=32'hFFFFFFFD;
// @7:74
  LUT4 \d_cnst_sn.un36_df  (
	.I0(inf_abs0_2[24]),
	.I1(inf_abs0_2[25]),
	.I2(inf_abs0_2[26]),
	.I3(inf_abs0_2[31]),
	.O(un36_df)
);
defparam \d_cnst_sn.un36_df .INIT=16'h0080;
// @7:105
  LUT5 \d_cnst_sn.m[0]  (
	.I0(datai[0]),
	.I1(inf_abs0_2[0]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(m_2[0])
);
defparam \d_cnst_sn.m[0] .INIT=32'hCACACACC;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_14_2135_a5_2  (
	.I0(datai[30]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.I5(g0_2_0_i2_lut6_2_O6),
	.O(N_3568)
);
defparam \d_cnst_sn.reg0_28_14_2135_a5_2 .INIT=64'h0000000000000008;
// @7:243
  LUT4 reg3_1_1_axb_31_cZ (
	.I0(datai[31]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(reg3_1_1_axb_31)
);
defparam reg3_1_1_axb_31_cZ.INIT=16'hDDDF;
// @7:97
  LUT6 \d_cnst_sn.r_4_3[29]  (
	.I0(reg0[29]),
	.I1(reg1[29]),
	.I2(reg2[29]),
	.I3(un3_reg3_cry_25),
	.I4(N_3_0),
	.I5(N_13),
	.O(r_4[29])
);
defparam \d_cnst_sn.r_4_3[29] .INIT=64'hF0F0AAAAFF00CCCC;
// @7:47
  LUT6_L \d_cnst_sn.N_36_i  (
	.I0(reg0[2]),
	.I1(reg1[2]),
	.I2(reg2[2]),
	.I3(reg3[2]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.LO(N_36_i)
);
defparam \d_cnst_sn.N_36_i .INIT=64'hFF00F0F0CCCCAAAA;
// @7:318
  LUT6 un11_reg0_axb_19_cZ (
	.I0(datai[19]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[19]),
	.O(un11_reg0_axb_19)
);
defparam un11_reg0_axb_19_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_18_cZ (
	.I0(datai[18]),
	.I1(inf_abs0_2[18]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[18]),
	.O(un11_reg0_axb_18)
);
defparam un11_reg0_axb_18_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_17_cZ (
	.I0(datai[17]),
	.I1(inf_abs0_2[17]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[17]),
	.O(un11_reg0_axb_17)
);
defparam un11_reg0_axb_17_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_16_cZ (
	.I0(datai[16]),
	.I1(inf_abs0_2[16]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[16]),
	.O(un11_reg0_axb_16)
);
defparam un11_reg0_axb_16_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_15_cZ (
	.I0(datai[15]),
	.I1(inf_abs0_2[15]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[15]),
	.O(un11_reg0_axb_15)
);
defparam un11_reg0_axb_15_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_14_cZ (
	.I0(datai[14]),
	.I1(inf_abs0_2[14]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[14]),
	.O(un11_reg0_axb_14)
);
defparam un11_reg0_axb_14_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_13_cZ (
	.I0(datai[13]),
	.I1(inf_abs0_2[13]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[13]),
	.O(un11_reg0_axb_13)
);
defparam un11_reg0_axb_13_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_12_cZ (
	.I0(datai[12]),
	.I1(inf_abs0_2[12]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[12]),
	.O(un11_reg0_axb_12)
);
defparam un11_reg0_axb_12_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_11_cZ (
	.I0(datai[11]),
	.I1(inf_abs0_2[11]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[11]),
	.O(un11_reg0_axb_11)
);
defparam un11_reg0_axb_11_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_10_cZ (
	.I0(datai[10]),
	.I1(inf_abs0_2[10]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[10]),
	.O(un11_reg0_axb_10)
);
defparam un11_reg0_axb_10_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_9_cZ (
	.I0(datai[9]),
	.I1(inf_abs0_2[9]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[9]),
	.O(un11_reg0_axb_9)
);
defparam un11_reg0_axb_9_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_8_cZ (
	.I0(datai[8]),
	.I1(inf_abs0_2[8]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[8]),
	.O(un11_reg0_axb_8)
);
defparam un11_reg0_axb_8_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_7_cZ (
	.I0(datai[7]),
	.I1(inf_abs0_2[7]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[7]),
	.O(un11_reg0_axb_7)
);
defparam un11_reg0_axb_7_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_6_cZ (
	.I0(datai[6]),
	.I1(inf_abs0_2[6]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[6]),
	.O(un11_reg0_axb_6)
);
defparam un11_reg0_axb_6_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_5_cZ (
	.I0(datai[5]),
	.I1(inf_abs0_2[5]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[5]),
	.O(un11_reg0_axb_5)
);
defparam un11_reg0_axb_5_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_4_cZ (
	.I0(datai[4]),
	.I1(inf_abs0_2[4]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[4]),
	.O(un11_reg0_axb_4)
);
defparam un11_reg0_axb_4_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_3_cZ (
	.I0(datai[3]),
	.I1(inf_abs0_2[3]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[3]),
	.O(un11_reg0_axb_3)
);
defparam un11_reg0_axb_3_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_2_cZ (
	.I0(datai[2]),
	.I1(inf_abs0_2[2]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(N_28),
	.O(un11_reg0_axb_2)
);
defparam un11_reg0_axb_2_cZ.INIT=64'h35353533CACACACC;
// @7:318
  LUT6 un11_reg0_axb_1_cZ (
	.I0(datai[1]),
	.I1(inf_abs0_2[1]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[1]),
	.O(un11_reg0_axb_1)
);
defparam un11_reg0_axb_1_cZ.INIT=64'h35353533CACACACC;
// @7:243
  LUT5 reg3_1_1_axb_19_cZ (
	.I0(datai[19]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_19)
);
defparam reg3_1_1_axb_19_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_18_cZ (
	.I0(datai[18]),
	.I1(inf_abs0_2[18]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_18)
);
defparam reg3_1_1_axb_18_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_17_cZ (
	.I0(datai[17]),
	.I1(inf_abs0_2[17]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_17)
);
defparam reg3_1_1_axb_17_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_16_cZ (
	.I0(datai[16]),
	.I1(inf_abs0_2[16]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_16)
);
defparam reg3_1_1_axb_16_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_15_cZ (
	.I0(datai[15]),
	.I1(inf_abs0_2[15]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_15)
);
defparam reg3_1_1_axb_15_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_14_cZ (
	.I0(datai[14]),
	.I1(inf_abs0_2[14]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_14)
);
defparam reg3_1_1_axb_14_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_13_cZ (
	.I0(datai[13]),
	.I1(inf_abs0_2[13]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_13)
);
defparam reg3_1_1_axb_13_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_12_cZ (
	.I0(datai[12]),
	.I1(inf_abs0_2[12]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_12)
);
defparam reg3_1_1_axb_12_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_11_cZ (
	.I0(datai[11]),
	.I1(inf_abs0_2[11]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_11)
);
defparam reg3_1_1_axb_11_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_10_cZ (
	.I0(datai[10]),
	.I1(inf_abs0_2[10]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_10)
);
defparam reg3_1_1_axb_10_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_9_cZ (
	.I0(datai[9]),
	.I1(inf_abs0_2[9]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_9)
);
defparam reg3_1_1_axb_9_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_8_cZ (
	.I0(datai[8]),
	.I1(inf_abs0_2[8]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_8)
);
defparam reg3_1_1_axb_8_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_7_cZ (
	.I0(datai[7]),
	.I1(inf_abs0_2[7]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_7)
);
defparam reg3_1_1_axb_7_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_6_cZ (
	.I0(datai[6]),
	.I1(inf_abs0_2[6]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_6)
);
defparam reg3_1_1_axb_6_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_5_cZ (
	.I0(datai[5]),
	.I1(inf_abs0_2[5]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_5)
);
defparam reg3_1_1_axb_5_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_4_cZ (
	.I0(datai[4]),
	.I1(inf_abs0_2[4]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_4)
);
defparam reg3_1_1_axb_4_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_3_cZ (
	.I0(datai[3]),
	.I1(inf_abs0_2[3]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_3)
);
defparam reg3_1_1_axb_3_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_2_cZ (
	.I0(datai[2]),
	.I1(inf_abs0_2[2]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_2)
);
defparam reg3_1_1_axb_2_cZ.INIT=32'h35353533;
// @7:243
  LUT5 reg3_1_1_axb_1_cZ (
	.I0(datai[1]),
	.I1(inf_abs0_2[1]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_1)
);
defparam reg3_1_1_axb_1_cZ.INIT=32'h35353533;
// @7:97
  LUT6 \d_cnst_sn.r_4_3[31]  (
	.I0(reg0[31]),
	.I1(reg1[31]),
	.I2(reg2[31]),
	.I3(inf_abs0_2[31]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.O(r_4[31])
);
defparam \d_cnst_sn.r_4_3[31] .INIT=64'hAA00AAF0AACCAAAA;
// @7:213
  LUT4 \d_cnst_sn.d_cnsts2  (
	.I0(inf_abs0_2[24]),
	.I1(inf_abs0_2[25]),
	.I2(inf_abs0_2[26]),
	.I3(inf_abs0_2[31]),
	.O(d_cnst_sm0)
);
defparam \d_cnst_sn.d_cnsts2 .INIT=16'h00BC;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_3_2492_0_cZ  (
	.I0(datai[19]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(N_3873_2),
	.I5(g0_2_0_i2_lut6_2_O6),
	.O(\d_cnst_sn.reg0_28_3_2492_0 )
);
defparam \d_cnst_sn.reg0_28_3_2492_0_cZ .INIT=64'h00CC000000A00000;
// @7:47
  LUT6 \d_cnst_sn.addr_20_iv_7_654_i_1_cZ  (
	.I0(reg1[0]),
	.I1(reg3[0]),
	.I2(state[0]),
	.I3(inf_abs0_2[0]),
	.I4(inf_abs0_2[27]),
	.I5(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_7_654_i_1 )
);
defparam \d_cnst_sn.addr_20_iv_7_654_i_1_cZ .INIT=64'h0303A35303F3A3F3;
// @7:212
  LUT5 \d_cnst_sn.reg3_4_sqmuxa_3_2  (
	.I0(inf_abs0_2[24]),
	.I1(inf_abs0_2[25]),
	.I2(inf_abs0_2[26]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg3_5_sqmuxa_2_1 )
);
defparam \d_cnst_sn.reg3_4_sqmuxa_3_2 .INIT=32'hFFFF007F;
// @7:74
  LUT5 \d_cnst_sn.reg2_16_11_a1[29]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[28]),
	.O(reg2_16_11_a1[29])
);
defparam \d_cnst_sn.reg2_16_11_a1[29] .INIT=32'h08000000;
// @7:103
  LUT6 \d_cnst_sn.b_cnst_0_x2  (
	.I0(N_3913),
	.I1(N_512_i),
	.I2(N_513_i),
	.I3(un11_r_cry[30]),
	.I4(un14_r_0_I_83),
	.I5(N_895),
	.O(N_3912)
);
defparam \d_cnst_sn.b_cnst_0_x2 .INIT=64'h5556595AA5A6A9AA;
// @7:318
  LUT6 un11_reg0_axb_0_cZ (
	.I0(datai[0]),
	.I1(inf_abs0_2[0]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.I5(r_4[0]),
	.O(un11_reg0_axb_0)
);
defparam un11_reg0_axb_0_cZ.INIT=64'h35353533CACACACC;
// @7:466
  LUT6 un3_t_axb_30_cZ (
	.I0(reg0[30]),
	.I1(reg1[30]),
	.I2(reg2[30]),
	.I3(inf_abs0_2[31]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.O(un3_t_axb_30)
);
defparam un3_t_axb_30_cZ.INIT=64'h55FF550F55335555;
// @7:466
  LUT6 un3_t_axb_29_cZ (
	.I0(reg0[29]),
	.I1(reg1[29]),
	.I2(reg2[29]),
	.I3(un3_reg3_cry_25),
	.I4(N_3_0),
	.I5(N_13),
	.O(un3_t_axb_29)
);
defparam un3_t_axb_29_cZ.INIT=64'h0F0F555500FF3333;
// @7:243
  LUT5 reg3_1_1_axb_0_cZ (
	.I0(datai[0]),
	.I1(inf_abs0_2[0]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.I4(inf_abs0_2[28]),
	.O(reg3_1_1_axb_0)
);
defparam reg3_1_1_axb_0_cZ.INIT=32'h35353533;
// @7:47
  LUT5 \d_cnst_sn.addr_4_sqmuxa_1_1  (
	.I0(inf_abs0_2[24]),
	.I1(inf_abs0_2[23]),
	.I2(inf_abs0_2[25]),
	.I3(inf_abs0_2[26]),
	.I4(inf_abs0_2[31]),
	.O(addr_4_sqmuxa_1_1)
);
defparam \d_cnst_sn.addr_4_sqmuxa_1_1 .INIT=32'h00002000;
// @7:466
  LUT6 \d_cnst_sn.r_4_i[31]  (
	.I0(reg0[31]),
	.I1(reg1[31]),
	.I2(reg2[31]),
	.I3(inf_abs0_2[31]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.O(r_4_i[31])
);
defparam \d_cnst_sn.r_4_i[31] .INIT=64'h55FF550F55335555;
// @7:466
  LUT6 un3_t_axb_31_cZ (
	.I0(reg0[31]),
	.I1(reg1[31]),
	.I2(reg2[31]),
	.I3(inf_abs0_2[31]),
	.I4(inf_abs0_2[29]),
	.I5(inf_abs0_2[30]),
	.O(un3_t_axb_31)
);
defparam un3_t_axb_31_cZ.INIT=64'h55FF550F55335555;
// @7:47
  LUT6 \d_cnst_sn.addr_20_iv_9_589_x2  (
	.I0(reg2[0]),
	.I1(reg1[0]),
	.I2(inf_abs0_2[0]),
	.I3(inf_abs0_2[31]),
	.I4(inf_abs0_2[27]),
	.I5(inf_abs0_2[28]),
	.O(N_2240_i)
);
defparam \d_cnst_sn.addr_20_iv_9_589_x2 .INIT=64'hF05AF03CF0F0F0F0;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_14_2135_1_a0_2_cZ  (
	.I0(b),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.I4(inf_abs0_2[27]),
	.I5(inf_abs0_2[28]),
	.O(\d_cnst_sn.reg0_28_14_2135_1_a0_2 )
);
defparam \d_cnst_sn.reg0_28_14_2135_1_a0_2_cZ .INIT=64'h00000000004000C0;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_0_cZ[25]  (
	.I0(N_512_i),
	.I1(N_513_i),
	.I2(N_514_i),
	.I3(m_2[25]),
	.I4(N_527_i),
	.I5(r_4[24]),
	.O(\d_cnst_sn.reg2_16_0 [25])
);
defparam \d_cnst_sn.reg2_16_0_cZ[25] .INIT=64'hFFFDFFFD3F3DFFFD;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_0_cZ[24]  (
	.I0(N_512_i),
	.I1(N_513_i),
	.I2(N_514_i),
	.I3(m_2[24]),
	.I4(N_527_i),
	.I5(r_4[23]),
	.O(\d_cnst_sn.reg2_16_0 [24])
);
defparam \d_cnst_sn.reg2_16_0_cZ[24] .INIT=64'hFFFDFFFD3F3DFFFD;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_0_cZ[23]  (
	.I0(N_512_i),
	.I1(N_513_i),
	.I2(N_514_i),
	.I3(m_2[23]),
	.I4(N_527_i),
	.I5(r_4[22]),
	.O(\d_cnst_sn.reg2_16_0 [23])
);
defparam \d_cnst_sn.reg2_16_0_cZ[23] .INIT=64'hFFFDFFFD3F3DFFFD;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_0_cZ[22]  (
	.I0(N_512_i),
	.I1(N_513_i),
	.I2(N_514_i),
	.I3(m_2[22]),
	.I4(N_527_i),
	.I5(r_4[21]),
	.O(\d_cnst_sn.reg2_16_0 [22])
);
defparam \d_cnst_sn.reg2_16_0_cZ[22] .INIT=64'hFFFDFFFD3F3DFFFD;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_0_cZ[21]  (
	.I0(N_512_i),
	.I1(N_513_i),
	.I2(N_514_i),
	.I3(m_2[21]),
	.I4(N_527_i),
	.I5(r_4[20]),
	.LO(\d_cnst_sn.reg2_16_0 [21])
);
defparam \d_cnst_sn.reg2_16_0_cZ[21] .INIT=64'hFFFDFFFD3F3DFFFD;
// @7:103
  LUT5 \d_cnst_sn.un1_b59  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.O(un1_b59)
);
defparam \d_cnst_sn.un1_b59 .INIT=32'h00000AC0;
// @7:103
  LUT5 \d_cnst_sn.un1_b57  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.O(un1_b57)
);
defparam \d_cnst_sn.un1_b57 .INIT=32'h00000530;
// @7:47
  LUT5 \d_cnst_sn.reg0_m9_i_a1  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[28]),
	.O(reg0_m9_i_a1)
);
defparam \d_cnst_sn.reg0_m9_i_a1 .INIT=32'h08000000;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a2[29]  (
	.I0(un3_reg3_cry_25),
	.I1(N_3913),
	.I2(N_512_i),
	.I3(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I4(m_2[29]),
	.I5(reg3_1_1[29]),
	.O(reg2_16_11_a2[29])
);
defparam \d_cnst_sn.reg2_16_11_a2[29] .INIT=64'hFE000E00F2000200;
// @7:47
  LUT6 \d_cnst_sn.addr_4_sqmuxa_1  (
	.I0(state[0]),
	.I1(inf_abs0_2[24]),
	.I2(inf_abs0_2[23]),
	.I3(inf_abs0_2[25]),
	.I4(inf_abs0_2[26]),
	.I5(inf_abs0_2[31]),
	.O(addr_4_sqmuxa_1)
);
defparam \d_cnst_sn.addr_4_sqmuxa_1 .INIT=64'h0000000008000000;
// @7:213
  LUT4 \d_cnst_sn.d_cnst_ss0  (
	.I0(inf_abs0_2[24]),
	.I1(inf_abs0_2[25]),
	.I2(inf_abs0_2[26]),
	.I3(inf_abs0_2[31]),
	.O(d_cnst[0])
);
defparam \d_cnst_sn.d_cnst_ss0 .INIT=16'h00BA;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_17_362_i_1_RNI7JD51  (
	.I0(inf_abs0_2[28]),
	.I1(un1_inf_abs0_10[10]),
	.I2(un1_inf_abs0_11[10]),
	.I3(N_2660_2),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I5(\d_cnst_sn.addr_20_iv_17_362_i_1 ),
	.LO(N_2119_i)
);
defparam \d_cnst_sn.addr_20_iv_17_362_i_1_RNI7JD51 .INIT=64'h00000000D0F0DDFF;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_16_389_i_1_RNIVH7K1  (
	.I0(inf_abs0_2[28]),
	.I1(un1_inf_abs0_10[9]),
	.I2(un1_inf_abs0_11[9]),
	.I3(N_2660_2),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I5(\d_cnst_sn.addr_20_iv_16_389_i_1 ),
	.LO(N_2139_i)
);
defparam \d_cnst_sn.addr_20_iv_16_389_i_1_RNIVH7K1 .INIT=64'h00000000D0F0DDFF;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_15_416_i_1_RNI9QLS1  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_inf_abs0_10[8]),
	.I4(un1_inf_abs0_11[8]),
	.I5(\d_cnst_sn.addr_20_iv_15_416_i_1 ),
	.LO(N_2159_i)
);
defparam \d_cnst_sn.addr_20_iv_15_416_i_1_RNI9QLS1 .INIT=64'h00000000FF7FDD5D;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_14_443_i_2_RNILKQI1  (
	.I0(reg3[7]),
	.I1(state[0]),
	.I2(inf_abs0_2[7]),
	.I3(inf_abs0_2[28]),
	.I4(\d_cnst_sn.addr_20_iv_14_443_i_2 ),
	.I5(N_2641),
	.LO(N_2179_i)
);
defparam \d_cnst_sn.addr_20_iv_14_443_i_2_RNILKQI1 .INIT=64'h000000000000EEE2;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_13_470_i_1_RNI3GLV1  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_inf_abs0_10[6]),
	.I4(un1_inf_abs0_11[6]),
	.I5(\d_cnst_sn.addr_20_iv_13_470_i_1 ),
	.LO(N_2199_i)
);
defparam \d_cnst_sn.addr_20_iv_13_470_i_1_RNI3GLV1 .INIT=64'h00000000FF7FDD5D;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_12_497_i_1_RNI9EOO1  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_inf_abs0_10[5]),
	.I4(un1_inf_abs0_11[5]),
	.I5(\d_cnst_sn.addr_20_iv_12_497_i_1 ),
	.LO(N_2219_i)
);
defparam \d_cnst_sn.addr_20_iv_12_497_i_1_RNI9EOO1 .INIT=64'h00000000FF7FDD5D;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_10_562_i_1_RNIS0IN1  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_inf_abs0_10[3]),
	.I4(un1_inf_abs0_11[3]),
	.I5(\d_cnst_sn.addr_20_iv_10_562_i_1 ),
	.LO(N_2267_i)
);
defparam \d_cnst_sn.addr_20_iv_10_562_i_1_RNIS0IN1 .INIT=64'h00000000FF7FDD5D;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_0_cZ[20]  (
	.I0(\d_cnst_sn.reg2_N_3_mux ),
	.I1(reg2_16_2_d[20]),
	.I2(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I3(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I4(r_4[19]),
	.I5(reg3_1_1[20]),
	.O(\d_cnst_sn.reg2_16_0 [20])
);
defparam \d_cnst_sn.reg2_16_0_cZ[20] .INIT=64'hEFEF00EF4F4F004F;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_10  (
	.I0(m_2[2]),
	.I1(m_2[1]),
	.I2(m_2[0]),
	.I3(r_4[0]),
	.I4(r_4[1]),
	.I5(N_28),
	.O(un14_r_0_N_70)
);
defparam \d_cnst_sn.un14_r_0_I_10 .INIT=64'h8008200240041001;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_42  (
	.I0(m_2[15]),
	.I1(m_2[16]),
	.I2(m_2[17]),
	.I3(r_4[15]),
	.I4(r_4[16]),
	.I5(r_4[17]),
	.O(un14_r_0_N_42)
);
defparam \d_cnst_sn.un14_r_0_I_42 .INIT=64'h8040201008040201;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_74  (
	.I0(m_2[3]),
	.I1(m_2[4]),
	.I2(m_2[5]),
	.I3(r_4[3]),
	.I4(r_4[4]),
	.I5(r_4[5]),
	.O(un14_r_0_N_14)
);
defparam \d_cnst_sn.un14_r_0_I_74 .INIT=64'h8040201008040201;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_34  (
	.I0(m_2[19]),
	.I1(m_2[20]),
	.I2(m_2[18]),
	.I3(r_4[19]),
	.I4(r_4[18]),
	.I5(r_4[20]),
	.O(un14_r_0_N_49)
);
defparam \d_cnst_sn.un14_r_0_I_34 .INIT=64'h8040080420100201;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_82  (
	.I0(m_2[12]),
	.I1(m_2[13]),
	.I2(m_2[14]),
	.I3(r_4[12]),
	.I4(r_4[13]),
	.I5(r_4[14]),
	.O(un14_r_0_N_7)
);
defparam \d_cnst_sn.un14_r_0_I_82 .INIT=64'h8040201008040201;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_58  (
	.I0(m_2[9]),
	.I1(m_2[10]),
	.I2(m_2[11]),
	.I3(r_4[11]),
	.I4(r_4[9]),
	.I5(r_4[10]),
	.O(un14_r_0_N_28)
);
defparam \d_cnst_sn.un14_r_0_I_58 .INIT=64'h8008400420021001;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_66  (
	.I0(m_2[7]),
	.I1(m_2[6]),
	.I2(m_2[8]),
	.I3(r_4[6]),
	.I4(r_4[8]),
	.I5(r_4[7]),
	.O(un14_r_0_N_21)
);
defparam \d_cnst_sn.un14_r_0_I_66 .INIT=64'h8020080240100401;
// @7:148
  LUT6 \d_cnst_sn.r_6[30]  (
	.I0(reg0[30]),
	.I1(reg1[30]),
	.I2(reg2[30]),
	.I3(N_3_0),
	.I4(r_4[31]),
	.I5(N_13),
	.O(r_6[30])
);
defparam \d_cnst_sn.r_6[30] .INIT=64'hF0AA000000CC0000;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_a1_1_lut6_2_RNIH32G2[7]  (
	.I0(N_3910),
	.I1(\d_cnst_sn.reg0_28_a0_1 [7]),
	.I2(m_2[7]),
	.I3(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I4(r_4[6]),
	.I5(reg3_1_1[7]),
	.O(\d_cnst_sn.reg0_1 [7])
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_RNIH32G2[7] .INIT=64'hF5F500F531310031;
// @7:128
  LUT6 \d_cnst_sn.un14_r_0_I_18  (
	.I0(m_2[29]),
	.I1(m_2[27]),
	.I2(m_2[28]),
	.I3(r_4[27]),
	.I4(r_4[28]),
	.I5(r_4[29]),
	.O(un14_r_0_N_63)
);
defparam \d_cnst_sn.un14_r_0_I_18 .INIT=64'h8020080240100401;
// @7:212
  LUT6 \d_cnst_sn.b_2_sqmuxa  (
	.I0(N_526_i),
	.I1(N_1901),
	.I2(N_513_i),
	.I3(N_514_i),
	.I4(un36_df),
	.I5(N_527_i),
	.O(b_2_sqmuxa)
);
defparam \d_cnst_sn.b_2_sqmuxa .INIT=64'h0000200000000000;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_18_335_i_1_RNI0IID1  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_inf_abs0_10[11]),
	.I4(un1_inf_abs0_11[11]),
	.I5(\d_cnst_sn.addr_20_iv_18_335_i_1 ),
	.LO(N_2099_i)
);
defparam \d_cnst_sn.addr_20_iv_18_335_i_1_RNI0IID1 .INIT=64'h00000000FF7FDD5D;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_6_863_i_0_lut6_2_RNI74TR  (
	.I0(\d_cnst_sn.addr_20_iv_6_863_i_0 ),
	.I1(un1_inf_abs0_10[19]),
	.I2(un1_inf_abs0_11[19]),
	.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),
	.I5(N_2641),
	.LO(N_2516_i)
);
defparam \d_cnst_sn.addr_20_iv_6_863_i_0_lut6_2_RNI74TR .INIT=64'h0000000040445055;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_1052_i_a6_2_0_lut6_2_RNIUHOV1  (
	.I0(\d_cnst_sn.addr_20_iv_5_890_i_0 ),
	.I1(un1_inf_abs0_10[18]),
	.I2(un1_inf_abs0_11[18]),
	.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),
	.I5(N_2641),
	.LO(N_2536_i)
);
defparam \d_cnst_sn.addr_20_iv_1052_i_a6_2_0_lut6_2_RNIUHOV1 .INIT=64'h0000000040445055;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_4_917_i_0_lut6_2_RNI13AS  (
	.I0(\d_cnst_sn.addr_20_iv_4_917_i_0 ),
	.I1(un1_inf_abs0_10[17]),
	.I2(un1_inf_abs0_11[17]),
	.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),
	.I5(N_2641),
	.LO(N_2556_i)
);
defparam \d_cnst_sn.addr_20_iv_4_917_i_0_lut6_2_RNI13AS .INIT=64'h0000000040445055;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_1052_i_a6_2_0_lut6_2_RNIMFOV1  (
	.I0(\d_cnst_sn.addr_20_iv_3_944_i_0 ),
	.I1(un1_inf_abs0_10[16]),
	.I2(un1_inf_abs0_11[16]),
	.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),
	.I5(N_2641),
	.LO(N_2576_i)
);
defparam \d_cnst_sn.addr_20_iv_1052_i_a6_2_0_lut6_2_RNIMFOV1 .INIT=64'h0000000040445055;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_2_971_i_0_lut6_2_RNIRAP31  (
	.I0(\d_cnst_sn.addr_20_iv_2_971_i_0 ),
	.I1(un1_inf_abs0_10[15]),
	.I2(un1_inf_abs0_11[15]),
	.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),
	.I5(N_2641),
	.LO(N_2596_i)
);
defparam \d_cnst_sn.addr_20_iv_2_971_i_0_lut6_2_RNIRAP31 .INIT=64'h0000000040445055;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_1_998_i_0_lut6_2_RNI11O41  (
	.I0(\d_cnst_sn.addr_20_iv_1_998_i_0 ),
	.I1(un1_inf_abs0_10[14]),
	.I2(un1_inf_abs0_11[14]),
	.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),
	.I5(N_2641),
	.LO(N_2616_i)
);
defparam \d_cnst_sn.addr_20_iv_1_998_i_0_lut6_2_RNI11O41 .INIT=64'h0000000040445055;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_0_1025_i_0_lut6_2_RNIS79S  (
	.I0(\d_cnst_sn.addr_20_iv_0_1025_i_0 ),
	.I1(un1_inf_abs0_10[13]),
	.I2(un1_inf_abs0_11[13]),
	.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),
	.I5(N_2641),
	.LO(N_2636_i)
);
defparam \d_cnst_sn.addr_20_iv_0_1025_i_0_lut6_2_RNIS79S .INIT=64'h0000000040445055;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_1052_i_0_lut6_2_RNIBHO61  (
	.I0(\d_cnst_sn.addr_20_iv_1052_i_0 ),
	.I1(un1_inf_abs0_10[12]),
	.I2(un1_inf_abs0_11[12]),
	.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),
	.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),
	.I5(N_2641),
	.LO(N_2656_i)
);
defparam \d_cnst_sn.addr_20_iv_1052_i_0_lut6_2_RNIBHO61 .INIT=64'h0000000040445055;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_0_1_0_cZ[28]  (
	.I0(\d_cnst_sn.reg2_16_0_1_tz [28]),
	.I1(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[27]),
	.I4(N_1363),
	.I5(un32_reg0_s_28),
	.O(\d_cnst_sn.reg2_16_0_1_0 [28])
);
defparam \d_cnst_sn.reg2_16_0_1_0_cZ[28] .INIT=64'hFF0F3303AA0A2202;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_0_1_0_cZ[27]  (
	.I0(\d_cnst_sn.reg2_16_0_1_tz [28]),
	.I1(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[26]),
	.I4(N_1362),
	.I5(un32_reg0_s_27),
	.O(\d_cnst_sn.reg2_16_0_1_0 [27])
);
defparam \d_cnst_sn.reg2_16_0_1_0_cZ[27] .INIT=64'hFF0F3303AA0A2202;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_0_1_0_cZ[26]  (
	.I0(\d_cnst_sn.reg2_16_0_1_tz [28]),
	.I1(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[25]),
	.I4(N_1361),
	.I5(un32_reg0_s_26),
	.O(\d_cnst_sn.reg2_16_0_1_0 [26])
);
defparam \d_cnst_sn.reg2_16_0_1_0_cZ[26] .INIT=64'hFF0F3303AA0A2202;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a3[17]  (
	.I0(N_3913),
	.I1(N_513_i),
	.I2(N_514_i),
	.I3(N_1352),
	.I4(un32_reg0_s_17),
	.I5(un11_reg0_s_17),
	.O(reg2_16_11_a3[17])
);
defparam \d_cnst_sn.reg2_16_11_a3[17] .INIT=64'h0003101320233033;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a3[19]  (
	.I0(N_3913),
	.I1(N_513_i),
	.I2(N_514_i),
	.I3(N_1354),
	.I4(un32_reg0_s_19),
	.I5(un11_reg0_s_19),
	.O(reg2_16_11_a3[19])
);
defparam \d_cnst_sn.reg2_16_11_a3[19] .INIT=64'h0003101320233033;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_11_a3[18]  (
	.I0(N_3913),
	.I1(N_513_i),
	.I2(N_514_i),
	.I3(N_1353),
	.I4(un32_reg0_s_18),
	.I5(un11_reg0_s_18),
	.O(reg2_16_11_a3[18])
);
defparam \d_cnst_sn.reg2_16_11_a3[18] .INIT=64'h0003101320233033;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[30]  (
	.I0(inf_abs0_2[22]),
	.I1(reg0_28_sn_m6_lut6_2_O5),
	.I2(N_513_i),
	.I3(N_527_i),
	.I4(N_1493),
	.I5(t_1[30]),
	.LO(reg2_16[30])
);
defparam \d_cnst_sn.reg2_16_11[30] .INIT=64'h0F0F00000F2F0020;
// @7:47
  LUT6 \d_cnst_sn.reg1_16_8_1837_0_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I3(m_2[27]),
	.I4(un32_reg0_s_27),
	.I5(un11_reg0_s_27),
	.O(\d_cnst_sn.reg1_16_8_1837_0 )
);
defparam \d_cnst_sn.reg1_16_8_1837_0_cZ .INIT=64'hFAAAF888F222F000;
// @7:47
  LUT6 \d_cnst_sn.reg1_16_7_1870_0_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I3(m_2[26]),
	.I4(un32_reg0_s_26),
	.I5(un11_reg0_s_26),
	.O(\d_cnst_sn.reg1_16_7_1870_0 )
);
defparam \d_cnst_sn.reg1_16_7_1870_0_cZ .INIT=64'hFAAAF888F222F000;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_9_2294_0_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I3(m_2[25]),
	.I4(un32_reg0_s_25),
	.I5(un11_reg0_s_25),
	.O(\d_cnst_sn.reg0_28_9_2294_0 )
);
defparam \d_cnst_sn.reg0_28_9_2294_0_cZ .INIT=64'hFAAAF888F222F000;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_7_2360_0_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I3(m_2[23]),
	.I4(un32_reg0_s_23),
	.I5(un11_reg0_s_23),
	.O(\d_cnst_sn.reg0_28_7_2360_0 )
);
defparam \d_cnst_sn.reg0_28_7_2360_0_cZ .INIT=64'hFAAAF888F222F000;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_6_2393_0_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I3(m_2[22]),
	.I4(un32_reg0_s_22),
	.I5(un11_reg0_s_22),
	.O(\d_cnst_sn.reg0_28_6_2393_0 )
);
defparam \d_cnst_sn.reg0_28_6_2393_0_cZ .INIT=64'hFAAAF888F222F000;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_5_2426_0_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I3(m_2[21]),
	.I4(un32_reg0_s_21),
	.I5(un11_reg0_s_21),
	.O(\d_cnst_sn.reg0_28_5_2426_0 )
);
defparam \d_cnst_sn.reg0_28_5_2426_0_cZ .INIT=64'hFAAAF888F222F000;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_8_2327_0_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I3(m_2[24]),
	.I4(un32_reg0_s_24),
	.I5(un11_reg0_s_24),
	.O(\d_cnst_sn.reg0_28_8_2327_0 )
);
defparam \d_cnst_sn.reg0_28_8_2327_0_cZ .INIT=64'hFAAAF888F222F000;
// @7:47
  LUT6 \d_cnst_sn.reg0_28_4_2459_0_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I3(m_2[20]),
	.I4(un32_reg0_s_20),
	.I5(un11_reg0_s_20),
	.O(\d_cnst_sn.reg0_28_4_2459_0 )
);
defparam \d_cnst_sn.reg0_28_4_2459_0_cZ .INIT=64'hFAAAF888F222F000;
// @7:47
  LUT5 \d_cnst_sn.reg0_28_3_2492_1_cZ  (
	.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),
	.I1(N_1033),
	.I2(\d_cnst_sn.reg0_28_3_2492_0 ),
	.I3(un32_reg0_s_19),
	.I4(un11_reg0_s_19),
	.O(\d_cnst_sn.reg0_28_3_2492_1 )
);
defparam \d_cnst_sn.reg0_28_3_2492_1_cZ .INIT=32'hFAF8F2F0;
// @7:74
  LUT6 \d_cnst_sn.reg2_16_1_0[29]  (
	.I0(N_512_i),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(reg2_16_11_a1[29]),
	.I3(reg2_16_11_a2[29]),
	.I4(un32_reg0_s_29),
	.I5(un11_reg0_s_29),
	.O(\d_cnst_sn.reg2_16_1 [29])
);
defparam \d_cnst_sn.reg2_16_1_0[29] .INIT=64'hFFFCFFF4FFF8FFF0;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[3]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1338),
	.I3(N_1370),
	.I4(N_1562),
	.I5(t_6[3]),
	.LO(reg2_16[3])
);
defparam \d_cnst_sn.reg2_16_11[3] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[4]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1339),
	.I3(N_1371),
	.I4(N_1563),
	.I5(t_6[4]),
	.LO(reg2_16[4])
);
defparam \d_cnst_sn.reg2_16_11[4] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[5]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1340),
	.I3(N_1372),
	.I4(N_1564),
	.I5(t_6[5]),
	.LO(reg2_16[5])
);
defparam \d_cnst_sn.reg2_16_11[5] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[6]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1341),
	.I3(N_1373),
	.I4(N_1565),
	.I5(t_6[6]),
	.LO(reg2_16[6])
);
defparam \d_cnst_sn.reg2_16_11[6] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[9]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1344),
	.I3(N_1376),
	.I4(N_1568),
	.I5(t_6[9]),
	.LO(reg2_16[9])
);
defparam \d_cnst_sn.reg2_16_11[9] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[10]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1345),
	.I3(N_1377),
	.I4(N_1569),
	.I5(t_6[10]),
	.LO(reg2_16[10])
);
defparam \d_cnst_sn.reg2_16_11[10] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[11]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1346),
	.I3(N_1378),
	.I4(N_1570),
	.I5(t_6[11]),
	.LO(reg2_16[11])
);
defparam \d_cnst_sn.reg2_16_11[11] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[12]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1347),
	.I3(N_1379),
	.I4(N_1571),
	.I5(t_6[12]),
	.LO(reg2_16[12])
);
defparam \d_cnst_sn.reg2_16_11[12] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[13]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1348),
	.I3(N_1380),
	.I4(N_1572),
	.I5(t_6[13]),
	.LO(reg2_16[13])
);
defparam \d_cnst_sn.reg2_16_11[13] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[14]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1349),
	.I3(N_1381),
	.I4(N_1573),
	.I5(t_6[14]),
	.LO(reg2_16[14])
);
defparam \d_cnst_sn.reg2_16_11[14] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[15]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1350),
	.I3(N_1382),
	.I4(N_1574),
	.I5(t_6[15]),
	.LO(reg2_16[15])
);
defparam \d_cnst_sn.reg2_16_11[15] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[16]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1351),
	.I3(N_1383),
	.I4(N_1575),
	.I5(t_6[16]),
	.LO(reg2_16[16])
);
defparam \d_cnst_sn.reg2_16_11[16] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.rd_18  (
	.I0(state[0]),
	.I1(N_7_i),
	.I2(N_513_i),
	.I3(N_514_i),
	.I4(un36_df),
	.I5(m7),
	.LO(rd_18)
);
defparam \d_cnst_sn.rd_18 .INIT=64'h55555555DDDDDFFF;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[8]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1343),
	.I3(N_1375),
	.I4(N_1567),
	.I5(t_6[8]),
	.LO(reg2_16[8])
);
defparam \d_cnst_sn.reg2_16_11[8] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[2]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1337),
	.I3(N_1369),
	.I4(N_1561),
	.I5(t_6[2]),
	.LO(reg2_16[2])
);
defparam \d_cnst_sn.reg2_16_11[2] .INIT=64'hFEBADC9876325410;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16_11[7]  (
	.I0(N_513_i),
	.I1(N_514_i),
	.I2(N_1342),
	.I3(N_1374),
	.I4(N_1566),
	.I5(t_6[7]),
	.LO(reg2_16[7])
);
defparam \d_cnst_sn.reg2_16_11[7] .INIT=64'hFEBADC9876325410;
// @7:47
  LUT6 \d_cnst_sn.addr_0_sqmuxa_1_i  (
	.I0(state[0]),
	.I1(N_7_i),
	.I2(N_513_i),
	.I3(N_514_i),
	.I4(un36_df),
	.I5(m7),
	.O(addr_0_sqmuxa_1_i)
);
defparam \d_cnst_sn.addr_0_sqmuxa_1_i .INIT=64'h77775555FFFFDFFF;
// @7:47
  LUT6 \d_cnst_sn.reg1_16_9_1804_3_tz_cZ  (
	.I0(\d_cnst_sn.reg0_28_12_2195_a6_1_2_0 ),
	.I1(\d_cnst_sn.reg0_m8_e_0 ),
	.I2(N_513_i),
	.I3(N_527_i),
	.I4(r_4[27]),
	.I5(reg3_1_1[28]),
	.O(\d_cnst_sn.reg1_16_9_1804_3_tz )
);
defparam \d_cnst_sn.reg1_16_9_1804_3_tz_cZ .INIT=64'hBBBBABBBB0B0A0B0;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[17]  (
	.I0(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(r_4[16]),
	.I3(t_1[17]),
	.I4(reg2_16_11_a2[17]),
	.I5(reg2_16_11_a3[17]),
	.LO(reg2_16[17])
);
defparam \d_cnst_sn.reg2_16[17] .INIT=64'h00000000000031F5;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[19]  (
	.I0(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(r_4[18]),
	.I3(t_1[19]),
	.I4(reg2_16_11_a2[19]),
	.I5(reg2_16_11_a3[19]),
	.LO(reg2_16[19])
);
defparam \d_cnst_sn.reg2_16[19] .INIT=64'h00000000000031F5;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[18]  (
	.I0(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(r_4[17]),
	.I3(t_1[18]),
	.I4(reg2_16_11_a2[18]),
	.I5(reg2_16_11_a3[18]),
	.LO(reg2_16[18])
);
defparam \d_cnst_sn.reg2_16[18] .INIT=64'h00000000000031F5;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[20]  (
	.I0(\d_cnst_sn.reg2_16_11_1_tz [28]),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(\d_cnst_sn.reg2_16_0 [20]),
	.I3(un11_reg0_s_20),
	.I4(\d_cnst_sn.reg2_16_1 [20]),
	.I5(t_1[20]),
	.LO(reg2_16[20])
);
defparam \d_cnst_sn.reg2_16[20] .INIT=64'h30200000F0A00000;
// @7:74
  LUT5_L \d_cnst_sn.reg2_16_0[28]  (
	.I0(\d_cnst_sn.reg2_16_11_1_tz [28]),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(un11_reg0_s_28),
	.I3(\d_cnst_sn.reg2_16_0_1_0 [28]),
	.I4(t_1[28]),
	.LO(reg2_16[28])
);
defparam \d_cnst_sn.reg2_16_0[28] .INIT=32'h3200FA00;
// @7:74
  LUT5_L \d_cnst_sn.reg2_16_0[27]  (
	.I0(\d_cnst_sn.reg2_16_11_1_tz [28]),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(un11_reg0_s_27),
	.I3(\d_cnst_sn.reg2_16_0_1_0 [27]),
	.I4(t_1[27]),
	.LO(reg2_16[27])
);
defparam \d_cnst_sn.reg2_16_0[27] .INIT=32'h3200FA00;
// @7:74
  LUT5_L \d_cnst_sn.reg2_16_0[26]  (
	.I0(\d_cnst_sn.reg2_16_11_1_tz [28]),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(un11_reg0_s_26),
	.I3(\d_cnst_sn.reg2_16_0_1_0 [26]),
	.I4(t_1[26]),
	.LO(reg2_16[26])
);
defparam \d_cnst_sn.reg2_16_0[26] .INIT=32'h3200FA00;
// @7:245
  LUT5_L \d_cnst_sn.un86_df  (
	.I0(d[0]),
	.I1(d[1]),
	.I2(un1_df_1),
	.I3(d_cnst[0]),
	.I4(d_cnst_sm0),
	.LO(un86_df)
);
defparam \d_cnst_sn.un86_df .INIT=32'h404F4040;
// @7:47
  LUT6_L \d_cnst_sn.reg0_28_4_2459  (
	.I0(\d_cnst_sn.reg0_28_2526_a5_1_0 ),
	.I1(\d_cnst_sn.reg1_16_8_1837_2_tz ),
	.I2(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I3(\d_cnst_sn.reg0_28_0 [20]),
	.I4(t_1[20]),
	.I5(\d_cnst_sn.reg0_28_4_2459_0 ),
	.LO(reg0_28_4_2459)
);
defparam \d_cnst_sn.reg0_28_4_2459 .INIT=64'hFFFFFFFF0E00EE00;
// @7:47
  LUT5_L \d_cnst_sn.reg1_16_8_1837  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_11_2228_a6_1_1 ),
	.I2(\d_cnst_sn.reg1_16_8_1837_3_1 ),
	.I3(t_1[27]),
	.I4(\d_cnst_sn.reg1_16_8_1837_0 ),
	.LO(reg1_16_8_1837)
);
defparam \d_cnst_sn.reg1_16_8_1837 .INIT=32'hFFFF54FC;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_7_2360  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_7_2360_3_1 ),
	.I2(\d_cnst_sn.reg0_28_7_2360_a6_1_1 ),
	.I3(t_1[23]),
	.I4(\d_cnst_sn.reg0_28_7_2360_0 ),
	.LO(reg0_28_7_2360)
);
defparam \d_cnst_sn.reg0_28_7_2360 .INIT=32'hFFFF54FC;
// @7:47
  LUT5_L \d_cnst_sn.reg1_16_7_1870  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_10_2261_a6_1_1 ),
	.I2(\d_cnst_sn.reg1_16_7_1870_3_1 ),
	.I3(t_1[26]),
	.I4(\d_cnst_sn.reg1_16_7_1870_0 ),
	.LO(reg1_16_7_1870)
);
defparam \d_cnst_sn.reg1_16_7_1870 .INIT=32'hFFFF54FC;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_5_2426  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_5_2426_3_1 ),
	.I2(\d_cnst_sn.reg0_28_5_2426_a6_1_1 ),
	.I3(t_1[21]),
	.I4(\d_cnst_sn.reg0_28_5_2426_0 ),
	.LO(reg0_28_5_2426)
);
defparam \d_cnst_sn.reg0_28_5_2426 .INIT=32'hFFFF54FC;
// @7:47
  LUT6_L \d_cnst_sn.reg0_28_3_2492  (
	.I0(\d_cnst_sn.reg0_28_2526_a5_1_0 ),
	.I1(\d_cnst_sn.reg1_16_8_1837_2_tz ),
	.I2(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I3(\d_cnst_sn.reg0_28_0 [19]),
	.I4(t_1[19]),
	.I5(\d_cnst_sn.reg0_28_3_2492_1 ),
	.LO(reg0_28_3_2492)
);
defparam \d_cnst_sn.reg0_28_3_2492 .INIT=64'hFFFFFFFF0E00EE00;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_6_2393  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_6_2393_3_1 ),
	.I2(\d_cnst_sn.reg0_28_6_2393_a6_1_1 ),
	.I3(t_1[22]),
	.I4(\d_cnst_sn.reg0_28_6_2393_0 ),
	.LO(reg0_28_6_2393)
);
defparam \d_cnst_sn.reg0_28_6_2393 .INIT=32'hFFFF54FC;
// @7:47
  LUT5_L \d_cnst_sn.reg0_28_9_2294  (
	.I0(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I1(\d_cnst_sn.reg0_28_9_2294_3_1 ),
	.I2(\d_cnst_sn.reg0_28_9_2294_a6_1_1 ),
	.I3(t_1[25]),
	.I4(\d_cnst_sn.reg0_28_9_2294_0 ),
	.LO(N_3673)
);
defparam \d_cnst_sn.reg0_28_9_2294 .INIT=32'hFFFF54FC;
// @7:47
  LUT6_L \d_cnst_sn.reg0_28_8_2327  (
	.I0(\d_cnst_sn.reg1_16_8_1837_2_tz ),
	.I1(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I2(reg0_28_7_d[24]),
	.I3(\d_cnst_sn.reg0_28_8_2327_a6_1_1 ),
	.I4(t_1[24]),
	.I5(\d_cnst_sn.reg0_28_8_2327_0 ),
	.LO(reg0_28_8_2327)
);
defparam \d_cnst_sn.reg0_28_8_2327 .INIT=64'hFFFFFFFF3320FFA8;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[29]  (
	.I0(\d_cnst_sn.reg0_m9_i_a0_0 ),
	.I1(N_514_i),
	.I2(N_527_i),
	.I3(t_1[29]),
	.I4(reg2_16_11_a3[29]),
	.I5(\d_cnst_sn.reg2_16_1 [29]),
	.LO(reg2_16[29])
);
defparam \d_cnst_sn.reg2_16[29] .INIT=64'hFFFFFFFFFFFF0008;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNI0TVT3_0[7]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg0_1 [7]),
	.I4(t_1[7]),
	.I5(N_1042),
	.LO(reg0_28[7])
);
defparam \d_cnst_sn.reg0_28_6_RNI0TVT3_0[7] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[25]  (
	.I0(\d_cnst_sn.b60_0 ),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(\d_cnst_sn.reg2_16_1 [25]),
	.I3(t_1[25]),
	.I4(reg2_16_11_a4[25]),
	.I5(N_1584),
	.LO(reg2_16[25])
);
defparam \d_cnst_sn.reg2_16[25] .INIT=64'h000030F000001050;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[24]  (
	.I0(\d_cnst_sn.b60_0 ),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(\d_cnst_sn.reg2_16_1 [24]),
	.I3(t_1[24]),
	.I4(reg2_16_11_a4[24]),
	.I5(N_1583),
	.LO(reg2_16[24])
);
defparam \d_cnst_sn.reg2_16[24] .INIT=64'h000030F000001050;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[23]  (
	.I0(\d_cnst_sn.b60_0 ),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(\d_cnst_sn.reg2_16_1 [23]),
	.I3(t_1[23]),
	.I4(reg2_16_11_a4[23]),
	.I5(N_1582),
	.LO(reg2_16[23])
);
defparam \d_cnst_sn.reg2_16[23] .INIT=64'h000030F000001050;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[22]  (
	.I0(\d_cnst_sn.b60_0 ),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(\d_cnst_sn.reg2_16_1 [22]),
	.I3(t_1[22]),
	.I4(reg2_16_11_a4[22]),
	.I5(N_1581),
	.LO(reg2_16[22])
);
defparam \d_cnst_sn.reg2_16[22] .INIT=64'h000030F000001050;
// @7:74
  LUT6_L \d_cnst_sn.reg2_16[21]  (
	.I0(\d_cnst_sn.b60_0 ),
	.I1(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I2(\d_cnst_sn.reg2_16_1 [21]),
	.I3(t_1[21]),
	.I4(reg2_16_11_a4[21]),
	.I5(N_1580),
	.LO(reg2_16[21])
);
defparam \d_cnst_sn.reg2_16[21] .INIT=64'h000030F000001050;
// @7:47
  LUT6_L b_e (
	.I0(b),
	.I1(state[0]),
	.I2(N_7_i),
	.I3(N_514_i),
	.I4(b_2_sqmuxa),
	.I5(N_3912),
	.LO(b_0)
);
defparam b_e.INIT=64'hA222AA2AE2E2EAEA;
// @7:103
  LUT6 \d_cnst_sn.un1_df_16_2  (
	.I0(d[0]),
	.I1(d[1]),
	.I2(un1_df_1),
	.I3(d_cnst[0]),
	.I4(d_cnst_sm0),
	.I5(un36_df),
	.O(un1_df_17_2)
);
defparam \d_cnst_sn.un1_df_16_2 .INIT=64'h000000008F808080;
  LUT6_L \d_cnst_sn.addr_4_sqmuxa_1_1_RNIB1022  (
	.I0(inf_abs0_2[4]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_inf_abs0_10[4]),
	.I4(un1_inf_abs0_11[4]),
	.I5(addr_4_sqmuxa_1_1),
	.LO(N_54)
);
defparam \d_cnst_sn.addr_4_sqmuxa_1_1_RNIB1022 .INIT=64'hFFFFFFFF04C435F5;
  LUT6_L \d_cnst_sn.addr_4_sqmuxa_1_1_RNI51022  (
	.I0(inf_abs0_2[2]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.I3(un1_inf_abs0_10[2]),
	.I4(un1_inf_abs0_11[2]),
	.I5(addr_4_sqmuxa_1_1),
	.LO(N_45)
);
defparam \d_cnst_sn.addr_4_sqmuxa_1_1_RNI51022 .INIT=64'hFFFFFFFF04C435F5;
// @7:169
  LUT6 \d_cnst_sn.reg0_28_a1_1_lut6_2_RNISV191_0[7]  (
	.I0(d[0]),
	.I1(d[1]),
	.I2(un1_df_1),
	.I3(N_3910),
	.I4(d_cnst[0]),
	.I5(d_cnst_sm0),
	.O(N_1132)
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_RNISV191_0[7] .INIT=64'h1000100010001F00;
// @7:169
  LUT6 \d_cnst_sn.reg0_28_a1_1_lut6_2_RNISV191[7]  (
	.I0(d[0]),
	.I1(d[1]),
	.I2(un1_df_1),
	.I3(N_3910),
	.I4(d_cnst[0]),
	.I5(d_cnst_sm0),
	.O(N_1270)
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_RNISV191[7] .INIT=64'h200020002F002000;
// @7:47
  LUT6_L \d_cnst_sn.reg1_16_9  (
	.I0(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),
	.I1(m_2[28]),
	.I2(\d_cnst_sn.reg0_28_7_a0_0 [9]),
	.I3(\d_cnst_sn.reg1_16_9_1804_3_tz ),
	.I4(t_1[28]),
	.I5(N_3614),
	.LO(reg1_16_9)
);
defparam \d_cnst_sn.reg1_16_9 .INIT=64'hFFFFFFFF8F88FF88;
// @7:92
  LUT6 \d_cnst_sn.reg3_1_sqmuxa  (
	.I0(N_7_i),
	.I1(N_1901),
	.I2(N_513_i),
	.I3(N_514_i),
	.I4(un36_df),
	.I5(un87_df),
	.O(reg3_1_sqmuxa)
);
defparam \d_cnst_sn.reg3_1_sqmuxa .INIT=64'h0000000100000000;
// @7:92
  LUT6 \d_cnst_sn.reg3_14_sqmuxa  (
	.I0(N_7_i),
	.I1(N_1901),
	.I2(N_513_i),
	.I3(N_514_i),
	.I4(un36_df),
	.I5(un87_df),
	.O(reg3_14_sqmuxa)
);
defparam \d_cnst_sn.reg3_14_sqmuxa .INIT=64'h0000100000000000;
// @7:47
  LUT6 \d_cnst_sn.un1_state_4_1_RNIH54E1  (
	.I0(d[0]),
	.I1(d[1]),
	.I2(un1_df_1),
	.I3(d_cnst[0]),
	.I4(d_cnst_sm0),
	.I5(\d_cnst_sn.un1_state_3_1 ),
	.O(un1_state_3_i)
);
defparam \d_cnst_sn.un1_state_4_1_RNIH54E1 .INIT=64'h0000000020202F20;
// @7:47
  LUT6 \d_cnst_sn.un1_state_4_1_RNIH54E1_0  (
	.I0(d[0]),
	.I1(d[1]),
	.I2(un1_df_1),
	.I3(d_cnst[0]),
	.I4(d_cnst_sm0),
	.I5(\d_cnst_sn.un1_state_3_1 ),
	.O(un1_state_4_i)
);
defparam \d_cnst_sn.un1_state_4_1_RNIH54E1_0 .INIT=64'h000000001010101F;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[15]  (
	.I0(m_2[15]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1050),
	.I4(N_1082),
	.LO(reg0_28[15])
);
defparam \d_cnst_sn.reg0_28[15] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[15]  (
	.I0(m_2[15]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1050),
	.I4(N_1082),
	.LO(reg1_16[15])
);
defparam \d_cnst_sn.reg1_16[15] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[1]  (
	.I0(m_2[1]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1036),
	.I4(N_1068),
	.LO(reg0_28[1])
);
defparam \d_cnst_sn.reg0_28[1] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[16]  (
	.I0(m_2[16]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1051),
	.I4(N_1083),
	.LO(reg0_28[16])
);
defparam \d_cnst_sn.reg0_28[16] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[18]  (
	.I0(m_2[18]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1053),
	.I4(N_1085),
	.LO(reg0_28[18])
);
defparam \d_cnst_sn.reg0_28[18] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[1]  (
	.I0(m_2[1]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1036),
	.I4(N_1068),
	.LO(reg1_16[1])
);
defparam \d_cnst_sn.reg1_16[1] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[16]  (
	.I0(m_2[16]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1051),
	.I4(N_1083),
	.LO(reg1_16[16])
);
defparam \d_cnst_sn.reg1_16[16] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[13]  (
	.I0(m_2[13]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1048),
	.I4(N_1080),
	.LO(reg0_28[13])
);
defparam \d_cnst_sn.reg0_28[13] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[13]  (
	.I0(m_2[13]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1048),
	.I4(N_1080),
	.LO(reg1_16[13])
);
defparam \d_cnst_sn.reg1_16[13] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[9]  (
	.I0(m_2[9]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1044),
	.I4(N_1076),
	.LO(reg0_28[9])
);
defparam \d_cnst_sn.reg0_28[9] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[10]  (
	.I0(m_2[10]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1045),
	.I4(N_1077),
	.LO(reg0_28[10])
);
defparam \d_cnst_sn.reg0_28[10] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[11]  (
	.I0(m_2[11]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1046),
	.I4(N_1078),
	.LO(reg0_28[11])
);
defparam \d_cnst_sn.reg0_28[11] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[12]  (
	.I0(m_2[12]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1047),
	.I4(N_1079),
	.LO(reg0_28[12])
);
defparam \d_cnst_sn.reg0_28[12] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg0_28[14]  (
	.I0(m_2[14]),
	.I1(N_3916),
	.I2(N_1132),
	.I3(N_1049),
	.I4(N_1081),
	.LO(reg0_28[14])
);
defparam \d_cnst_sn.reg0_28[14] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[2]  (
	.I0(m_2[2]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1037),
	.I4(N_1069),
	.LO(reg1_16[2])
);
defparam \d_cnst_sn.reg1_16[2] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[9]  (
	.I0(m_2[9]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1044),
	.I4(N_1076),
	.LO(reg1_16[9])
);
defparam \d_cnst_sn.reg1_16[9] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[10]  (
	.I0(m_2[10]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1045),
	.I4(N_1077),
	.LO(reg1_16[10])
);
defparam \d_cnst_sn.reg1_16[10] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[11]  (
	.I0(m_2[11]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1046),
	.I4(N_1078),
	.LO(reg1_16[11])
);
defparam \d_cnst_sn.reg1_16[11] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[12]  (
	.I0(m_2[12]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1047),
	.I4(N_1079),
	.LO(reg1_16[12])
);
defparam \d_cnst_sn.reg1_16[12] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[14]  (
	.I0(m_2[14]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1049),
	.I4(N_1081),
	.LO(reg1_16[14])
);
defparam \d_cnst_sn.reg1_16[14] .INIT=32'hAFA3ACA0;
// @7:74
  LUT5_L \d_cnst_sn.reg1_16[17]  (
	.I0(m_2[17]),
	.I1(N_3916),
	.I2(N_1270),
	.I3(N_1052),
	.I4(N_1084),
	.LO(reg1_16[17])
);
defparam \d_cnst_sn.reg1_16[17] .INIT=32'hAFA3ACA0;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_a0_0[21]  (
	.I0(N_7_i),
	.I1(N_1901),
	.I2(N_513_i),
	.I3(N_514_i),
	.I4(un1_df_17_2),
	.I5(rd_4_sqmuxa),
	.O(reg3_17_sn_N_5)
);
defparam \d_cnst_sn.reg3_17_a0_0[21] .INIT=64'h00000000EFFFFFFF;
// @7:47
  LUT6 \d_cnst_sn.un86_df_RNIN5BD2  (
	.I0(state[0]),
	.I1(N_7_i),
	.I2(N_1892),
	.I3(un36_df),
	.I4(N_1890),
	.I5(un86_df),
	.O(un1_state_1_0_i)
);
defparam \d_cnst_sn.un86_df_RNIN5BD2 .INIT=64'h0002000200000002;
// @7:103
  LUT3 \d_cnst_sn.reg3_17_1[1]  (
	.I0(reg3[1]),
	.I1(reg3_1_1[1]),
	.I2(reg3_1_sqmuxa),
	.O(N_1689)
);
defparam \d_cnst_sn.reg3_17_1[1] .INIT=8'hCA;
// @7:103
  LUT3 \d_cnst_sn.reg3_17_1[2]  (
	.I0(reg3[2]),
	.I1(reg3_1_1[2]),
	.I2(reg3_1_sqmuxa),
	.O(N_1690)
);
defparam \d_cnst_sn.reg3_17_1[2] .INIT=8'hCA;
// @7:103
  LUT3 \d_cnst_sn.reg3_17_1[0]  (
	.I0(reg3[0]),
	.I1(m_2[0]),
	.I2(reg3_1_sqmuxa),
	.O(N_1688)
);
defparam \d_cnst_sn.reg3_17_1[0] .INIT=8'hCA;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_7_a1_RNIGOF53[18]  (
	.I0(N_513_i),
	.I1(m_2[18]),
	.I2(N_3916),
	.I3(reg0_28_7_a1[18]),
	.I4(N_1270),
	.I5(reg3_1_1[18]),
	.O(\d_cnst_sn.reg1_0 [18])
);
defparam \d_cnst_sn.reg0_28_7_a1_RNIGOF53[18] .INIT=64'hCCCCF0FFCCCCF0FA;
// @7:74
  LUT6 \d_cnst_sn.reg0_28_7_a1_RNIDMF53[17]  (
	.I0(N_513_i),
	.I1(m_2[17]),
	.I2(N_3916),
	.I3(reg0_28_7_a1[17]),
	.I4(N_1132),
	.I5(reg3_1_1[17]),
	.O(\d_cnst_sn.reg0_0 [17])
);
defparam \d_cnst_sn.reg0_28_7_a1_RNIDMF53[17] .INIT=64'hCCCCF0FFCCCCF0FA;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNI3QJL3[8]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[8]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[7]),
	.I4(reg3_1_1[8]),
	.I5(N_1132),
	.O(\d_cnst_sn.reg0_1 [8])
);
defparam \d_cnst_sn.m_2_RNI3QJL3[8] .INIT=64'hCCCCCCCCFF0F5505;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNI3QJL3_0[8]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[8]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[7]),
	.I4(reg3_1_1[8]),
	.I5(N_1270),
	.O(\d_cnst_sn.reg1_1 [8])
);
defparam \d_cnst_sn.m_2_RNI3QJL3_0[8] .INIT=64'hCCCCCCCCFF0F5505;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNIPHJL3[6]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[6]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[5]),
	.I4(reg3_1_1[6]),
	.I5(N_1132),
	.O(\d_cnst_sn.reg0_1 [6])
);
defparam \d_cnst_sn.m_2_RNIPHJL3[6] .INIT=64'hCCCCCCCCFF0F5505;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNIPHJL3_0[6]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[6]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[5]),
	.I4(reg3_1_1[6]),
	.I5(N_1270),
	.O(\d_cnst_sn.reg1_1 [6])
);
defparam \d_cnst_sn.m_2_RNIPHJL3_0[6] .INIT=64'hCCCCCCCCFF0F5505;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNIGF2R3[5]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[5]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[4]),
	.I4(reg3_1_1[5]),
	.I5(N_1132),
	.O(\d_cnst_sn.reg0_1 [5])
);
defparam \d_cnst_sn.m_2_RNIGF2R3[5] .INIT=64'hCCCCCCCCFF0F5505;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNIGF2R3_0[5]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[5]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[4]),
	.I4(reg3_1_1[5]),
	.I5(N_1270),
	.O(\d_cnst_sn.reg1_1 [5])
);
defparam \d_cnst_sn.m_2_RNIGF2R3_0[5] .INIT=64'hCCCCCCCCFF0F5505;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNI0T1N3[4]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[4]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[3]),
	.I4(reg3_1_1[4]),
	.I5(N_1270),
	.O(\d_cnst_sn.reg1_1 [4])
);
defparam \d_cnst_sn.m_2_RNI0T1N3[4] .INIT=64'hCCCCCCCCFF0F5505;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNI0T1N3_0[4]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[4]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(r_4[3]),
	.I4(reg3_1_1[4]),
	.I5(N_1132),
	.O(\d_cnst_sn.reg0_1 [4])
);
defparam \d_cnst_sn.m_2_RNI0T1N3_0[4] .INIT=64'hCCCCCCCCFF0F5505;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNIV5355[3]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[3]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(reg3_1_1[3]),
	.I4(N_28),
	.I5(N_1270),
	.O(\d_cnst_sn.reg1_1 [3])
);
defparam \d_cnst_sn.m_2_RNIV5355[3] .INIT=64'hCCCCCCCCFF550F05;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNIV5355_0[3]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[3]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(reg3_1_1[3]),
	.I4(N_28),
	.I5(N_1132),
	.O(\d_cnst_sn.reg0_1 [3])
);
defparam \d_cnst_sn.m_2_RNIV5355_0[3] .INIT=64'hCCCCCCCCFF550F05;
// @7:74
  LUT6 \d_cnst_sn.m_2_RNIMK1N3[2]  (
	.I0(\d_cnst_sn.reg1_16_a2_0 [5]),
	.I1(m_2[2]),
	.I2(\d_cnst_sn.reg0_28_a1_1 [4]),
	.I3(reg3_1_1[2]),
	.I4(r_4[1]),
	.I5(N_1132),
	.O(\d_cnst_sn.reg0_1 [2])
);
defparam \d_cnst_sn.m_2_RNIMK1N3[2] .INIT=64'hCCCCCCCCFF550F05;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_9_589_x2_RNIPBNN3  (
	.I0(reg3[4]),
	.I1(state[0]),
	.I2(inf_abs0_2[31]),
	.I3(N_2240_i),
	.I4(addr_4_sqmuxa_1_1),
	.I5(N_54),
	.LO(N_56_i)
);
defparam \d_cnst_sn.addr_20_iv_9_589_x2_RNIPBNN3 .INIT=64'hEE22E222EEEEEEEE;
// @7:47
  LUT6_L \d_cnst_sn.addr_20_iv_9_589_x2_RNIH9NN3  (
	.I0(reg3[2]),
	.I1(state[0]),
	.I2(inf_abs0_2[31]),
	.I3(N_2240_i),
	.I4(addr_4_sqmuxa_1_1),
	.I5(N_45),
	.LO(N_47_i)
);
defparam \d_cnst_sn.addr_20_iv_9_589_x2_RNIH9NN3 .INIT=64'hEE22E222EEEEEEEE;
// @7:103
  LUT5 \d_cnst_sn.reg3_N_7_i_RNO  (
	.I0(reg3[3]),
	.I1(inf_abs0_2[3]),
	.I2(reg3_1_1[3]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_N_7_i_RNO)
);
defparam \d_cnst_sn.reg3_N_7_i_RNO .INIT=32'h330F33AA;
// @7:103
  LUT5 \d_cnst_sn.reg3_1_sqmuxa_RNIEMUH1  (
	.I0(un3_reg3_s_1),
	.I1(inf_abs0_2[4]),
	.I2(reg3_1_1[4]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_1_sqmuxa_RNIEMUH1)
);
defparam \d_cnst_sn.reg3_1_sqmuxa_RNIEMUH1 .INIT=32'h330F3355;
// @7:103
  LUT5 \d_cnst_sn.reg3_1_sqmuxa_RNIHMUH1  (
	.I0(un3_reg3_s_2),
	.I1(inf_abs0_2[5]),
	.I2(reg3_1_1[5]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_1_sqmuxa_RNIHMUH1)
);
defparam \d_cnst_sn.reg3_1_sqmuxa_RNIHMUH1 .INIT=32'h330F3355;
// @7:103
  LUT5 \d_cnst_sn.reg3_1_sqmuxa_RNINMUH1  (
	.I0(un3_reg3_s_4),
	.I1(inf_abs0_2[7]),
	.I2(reg3_1_1[7]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_1_sqmuxa_RNINMUH1)
);
defparam \d_cnst_sn.reg3_1_sqmuxa_RNINMUH1 .INIT=32'h330F3355;
// @7:103
  LUT5 \d_cnst_sn.reg3_1_sqmuxa_RNIKMUH1  (
	.I0(un3_reg3_s_3),
	.I1(inf_abs0_2[6]),
	.I2(reg3_1_1[6]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_1_sqmuxa_RNIKMUH1)
);
defparam \d_cnst_sn.reg3_1_sqmuxa_RNIKMUH1 .INIT=32'h330F3355;
// @7:103
  LUT5 \d_cnst_sn.reg3_1_sqmuxa_RNITMUH1  (
	.I0(un3_reg3_s_6),
	.I1(inf_abs0_2[9]),
	.I2(reg3_1_1[9]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_1_sqmuxa_RNITMUH1)
);
defparam \d_cnst_sn.reg3_1_sqmuxa_RNITMUH1 .INIT=32'h330F3355;
// @7:103
  LUT5 \d_cnst_sn.reg3_1_sqmuxa_RNIQMUH1  (
	.I0(un3_reg3_s_5),
	.I1(inf_abs0_2[8]),
	.I2(reg3_1_1[8]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_1_sqmuxa_RNIQMUH1)
);
defparam \d_cnst_sn.reg3_1_sqmuxa_RNIQMUH1 .INIT=32'h330F3355;
// @7:103
  LUT5 \d_cnst_sn.reg3_1_sqmuxa_RNIE1DM1  (
	.I0(un3_reg3_s_7),
	.I1(inf_abs0_2[10]),
	.I2(reg3_1_1[10]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_1_sqmuxa_RNIE1DM1)
);
defparam \d_cnst_sn.reg3_1_sqmuxa_RNIE1DM1 .INIT=32'h330F3355;
// @7:103
  LUT5 \d_cnst_sn.reg3_1_sqmuxa_RNIH1DM1  (
	.I0(un3_reg3_s_8),
	.I1(inf_abs0_2[11]),
	.I2(reg3_1_1[11]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.O(reg3_1_sqmuxa_RNIH1DM1)
);
defparam \d_cnst_sn.reg3_1_sqmuxa_RNIH1DM1 .INIT=32'h330F3355;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[1]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(un11_reg0_s_1),
	.I3(un32_reg0_s_1),
	.I4(N_1658),
	.LO(N_1813)
);
defparam \d_cnst_sn.reg3_17_5[1] .INIT=32'hFEDC3210;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[27]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1684),
	.I3(un32_reg0_s_27),
	.I4(un11_reg0_s_27),
	.LO(N_1839)
);
defparam \d_cnst_sn.reg3_17_5[27] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[28]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1685),
	.I3(un32_reg0_s_28),
	.I4(un11_reg0_s_28),
	.LO(N_1840)
);
defparam \d_cnst_sn.reg3_17_5[28] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[16]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1673),
	.I3(un32_reg0_s_16),
	.I4(un11_reg0_s_16),
	.LO(N_1828)
);
defparam \d_cnst_sn.reg3_17_5[16] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[9]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1666),
	.I3(un32_reg0_s_9),
	.I4(un11_reg0_s_9),
	.O(N_1821)
);
defparam \d_cnst_sn.reg3_17_5[9] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[19]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1676),
	.I3(un32_reg0_s_19),
	.I4(un11_reg0_s_19),
	.LO(N_1831)
);
defparam \d_cnst_sn.reg3_17_5[19] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[20]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1677),
	.I3(un32_reg0_s_20),
	.I4(un11_reg0_s_20),
	.LO(N_1832)
);
defparam \d_cnst_sn.reg3_17_5[20] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[14]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1671),
	.I3(un32_reg0_s_14),
	.I4(un11_reg0_s_14),
	.LO(N_1826)
);
defparam \d_cnst_sn.reg3_17_5[14] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[18]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1675),
	.I3(un32_reg0_s_18),
	.I4(un11_reg0_s_18),
	.LO(N_1830)
);
defparam \d_cnst_sn.reg3_17_5[18] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[5]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1662),
	.I3(un32_reg0_s_5),
	.I4(un11_reg0_s_5),
	.O(N_1817)
);
defparam \d_cnst_sn.reg3_17_5[5] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[12]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1669),
	.I3(un32_reg0_s_12),
	.I4(un11_reg0_s_12),
	.LO(N_1824)
);
defparam \d_cnst_sn.reg3_17_5[12] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[17]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1674),
	.I3(un32_reg0_s_17),
	.I4(un11_reg0_s_17),
	.LO(N_1829)
);
defparam \d_cnst_sn.reg3_17_5[17] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[10]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1667),
	.I3(un32_reg0_s_10),
	.I4(un11_reg0_s_10),
	.O(N_1822)
);
defparam \d_cnst_sn.reg3_17_5[10] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[11]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1668),
	.I3(un32_reg0_s_11),
	.I4(un11_reg0_s_11),
	.O(N_1823)
);
defparam \d_cnst_sn.reg3_17_5[11] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[2]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(un11_reg0_s_2),
	.I3(un32_reg0_s_2),
	.I4(N_1659),
	.LO(N_1814)
);
defparam \d_cnst_sn.reg3_17_5[2] .INIT=32'hFEDC3210;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[6]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1663),
	.I3(un32_reg0_s_6),
	.I4(un11_reg0_s_6),
	.O(N_1818)
);
defparam \d_cnst_sn.reg3_17_5[6] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[8]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1665),
	.I3(un32_reg0_s_8),
	.I4(un11_reg0_s_8),
	.O(N_1820)
);
defparam \d_cnst_sn.reg3_17_5[8] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[3]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(un32_reg0_s_3),
	.I3(un11_reg0_s_3),
	.I4(N_1660),
	.O(N_1815)
);
defparam \d_cnst_sn.reg3_17_5[3] .INIT=32'hFDEC3120;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[15]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1672),
	.I3(un32_reg0_s_15),
	.I4(un11_reg0_s_15),
	.LO(N_1827)
);
defparam \d_cnst_sn.reg3_17_5[15] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[26]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1683),
	.I3(un32_reg0_s_26),
	.I4(un11_reg0_s_26),
	.LO(N_1838)
);
defparam \d_cnst_sn.reg3_17_5[26] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17_5[25]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1682),
	.I3(un32_reg0_s_25),
	.I4(un11_reg0_s_25),
	.LO(N_1837)
);
defparam \d_cnst_sn.reg3_17_5[25] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[7]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1664),
	.I3(un32_reg0_s_7),
	.I4(un11_reg0_s_7),
	.O(N_1819)
);
defparam \d_cnst_sn.reg3_17_5[7] .INIT=32'hF3D1E2C0;
// @7:103
  LUT5 \d_cnst_sn.reg3_17_5[4]  (
	.I0(un1_df_16),
	.I1(N_1810),
	.I2(N_1661),
	.I3(un32_reg0_s_4),
	.I4(un11_reg0_s_4),
	.O(N_1816)
);
defparam \d_cnst_sn.reg3_17_5[4] .INIT=32'hF3D1E2C0;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_0_cZ[28]  (
	.I0(un3_reg3_s_25),
	.I1(\d_cnst_sn.reg3_17_4_a2_0 [28]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_1[28]),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_14_sqmuxa),
	.O(\d_cnst_sn.reg3_17_6_0 [28])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[28] .INIT=64'hCCCCCCCC0F000A0A;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_0_cZ[27]  (
	.I0(un3_reg3_s_24),
	.I1(\d_cnst_sn.reg3_17_4_a2_0 [27]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_1[27]),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_14_sqmuxa),
	.O(\d_cnst_sn.reg3_17_6_0 [27])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[27] .INIT=64'hCCCCCCCC0F000A0A;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_1_cZ[18]  (
	.I0(un3_reg3_s_15),
	.I1(reg3_1_1[18]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.I5(\d_cnst_sn.reg3_17_6_0 [18]),
	.O(\d_cnst_sn.reg3_17_6_1 [18])
);
defparam \d_cnst_sn.reg3_17_6_1_cZ[18] .INIT=64'hFFFFFCFA00000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_1_cZ[19]  (
	.I0(un3_reg3_s_16),
	.I1(reg3_1_1[19]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.I5(\d_cnst_sn.reg3_17_6_0 [19]),
	.O(\d_cnst_sn.reg3_17_6_1 [19])
);
defparam \d_cnst_sn.reg3_17_6_1_cZ[19] .INIT=64'hFFFFFCFA00000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_0_cZ[26]  (
	.I0(un3_reg3_s_23),
	.I1(\d_cnst_sn.reg3_17_4_a2_0 [26]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_1[26]),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_14_sqmuxa),
	.O(\d_cnst_sn.reg3_17_6_0 [26])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[26] .INIT=64'hCCCCCCCC0F000A0A;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_1_cZ[17]  (
	.I0(un3_reg3_s_14),
	.I1(reg3_1_1[17]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.I5(\d_cnst_sn.reg3_17_6_0 [17]),
	.O(\d_cnst_sn.reg3_17_6_1 [17])
);
defparam \d_cnst_sn.reg3_17_6_1_cZ[17] .INIT=64'hFFFFFCFA00000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_0_cZ[25]  (
	.I0(un3_reg3_s_22),
	.I1(\d_cnst_sn.reg3_17_4_a2_0 [25]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_1[25]),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_14_sqmuxa),
	.O(\d_cnst_sn.reg3_17_6_0 [25])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[25] .INIT=64'hCCCCCCCC0F000A0A;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_1_cZ[16]  (
	.I0(un3_reg3_s_13),
	.I1(reg3_1_1[16]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.I5(\d_cnst_sn.reg3_17_6_0 [16]),
	.O(\d_cnst_sn.reg3_17_6_1 [16])
);
defparam \d_cnst_sn.reg3_17_6_1_cZ[16] .INIT=64'hFFFFFCFA00000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_1_cZ[15]  (
	.I0(un3_reg3_s_12),
	.I1(reg3_1_1[15]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.I5(\d_cnst_sn.reg3_17_6_0 [15]),
	.O(\d_cnst_sn.reg3_17_6_1 [15])
);
defparam \d_cnst_sn.reg3_17_6_1_cZ[15] .INIT=64'hFFFFFCFA00000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_1_cZ[14]  (
	.I0(un3_reg3_s_11),
	.I1(reg3_1_1[14]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.I5(\d_cnst_sn.reg3_17_6_0 [14]),
	.O(\d_cnst_sn.reg3_17_6_1 [14])
);
defparam \d_cnst_sn.reg3_17_6_1_cZ[14] .INIT=64'hFFFFFCFA00000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_1_cZ[13]  (
	.I0(un3_reg3_s_10),
	.I1(reg3_1_1[13]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.I5(\d_cnst_sn.reg3_17_6_0 [13]),
	.O(\d_cnst_sn.reg3_17_6_1 [13])
);
defparam \d_cnst_sn.reg3_17_6_1_cZ[13] .INIT=64'hFFFFFCFA00000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_0_cZ[20]  (
	.I0(un3_reg3_s_17),
	.I1(\d_cnst_sn.reg3_17_4_a2_0 [20]),
	.I2(reg3_1_1[20]),
	.I3(rd_4_sqmuxa),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_14_sqmuxa),
	.O(\d_cnst_sn.reg3_17_6_0 [20])
);
defparam \d_cnst_sn.reg3_17_6_0_cZ[20] .INIT=64'hCCCCCCCC00F000AA;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_6_1_cZ[12]  (
	.I0(un3_reg3_s_9),
	.I1(reg3_1_1[12]),
	.I2(rd_4_sqmuxa),
	.I3(reg3_1_sqmuxa),
	.I4(reg3_14_sqmuxa),
	.I5(\d_cnst_sn.reg3_17_6_0 [12]),
	.O(\d_cnst_sn.reg3_17_6_1 [12])
);
defparam \d_cnst_sn.reg3_17_6_1_cZ[12] .INIT=64'hFFFFFCFA00000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_a0[24]  (
	.I0(un3_reg3_s_21),
	.I1(reg3_1_1[24]),
	.I2(N_1810),
	.I3(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_17_sn_N_5),
	.O(reg3_17_a0[24])
);
defparam \d_cnst_sn.reg3_17_a0[24] .INIT=64'hC000A00000000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_a0[23]  (
	.I0(un3_reg3_s_20),
	.I1(reg3_1_1[23]),
	.I2(N_1810),
	.I3(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_17_sn_N_5),
	.O(reg3_17_a0[23])
);
defparam \d_cnst_sn.reg3_17_a0[23] .INIT=64'hC000A00000000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_a0[22]  (
	.I0(un3_reg3_s_19),
	.I1(reg3_1_1[22]),
	.I2(N_1810),
	.I3(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_17_sn_N_5),
	.O(reg3_17_a0[22])
);
defparam \d_cnst_sn.reg3_17_a0[22] .INIT=64'hC000A00000000000;
// @7:103
  LUT6 \d_cnst_sn.reg3_17_a0[21]  (
	.I0(un3_reg3_s_18),
	.I1(reg3_1_1[21]),
	.I2(N_1810),
	.I3(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I4(reg3_1_sqmuxa),
	.I5(reg3_17_sn_N_5),
	.O(reg3_17_a0[21])
);
defparam \d_cnst_sn.reg3_17_a0[21] .INIT=64'hC000A00000000000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[1]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_17_sn_N_5),
	.I3(N_1689),
	.I4(N_1751),
	.I5(N_1813),
	.LO(reg3_17[1])
);
defparam \d_cnst_sn.reg3_17[1] .INIT=64'hFF7FF77788088000;
// @7:103
  LUT5_L \d_cnst_sn.reg3_17[2]  (
	.I0(reg3_17_sn_N_5),
	.I1(N_1690),
	.I2(N_1841),
	.I3(N_1752),
	.I4(N_1814),
	.LO(reg3_17[2])
);
defparam \d_cnst_sn.reg3_17[2] .INIT=32'hDF8FD080;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[0]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_17_sn_N_5),
	.I3(N_1812),
	.I4(N_1688),
	.I5(N_1750),
	.LO(reg3_17[0])
);
defparam \d_cnst_sn.reg3_17[0] .INIT=64'hFF887F08F7807700;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNI6R0J6_0[3]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg0_1 [3]),
	.I4(t_1[3]),
	.I5(N_1038),
	.LO(reg0_28[3])
);
defparam \d_cnst_sn.reg0_28_6_RNI6R0J6_0[3] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNIR8V45[2]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg0_1 [2]),
	.I4(t_1[2]),
	.I5(N_1037),
	.LO(reg0_28[2])
);
defparam \d_cnst_sn.reg0_28_6_RNIR8V45[2] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNI6R0J6[3]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg1_1 [3]),
	.I4(t_1[3]),
	.I5(N_1038),
	.LO(reg1_16[3])
);
defparam \d_cnst_sn.reg0_28_6_RNI6R0J6[3] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNIKKH35[8]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg0_1 [8]),
	.I4(t_1[8]),
	.I5(N_1043),
	.LO(reg0_28[8])
);
defparam \d_cnst_sn.reg0_28_6_RNIKKH35[8] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNIKKH35_0[8]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg1_1 [8]),
	.I4(t_1[8]),
	.I5(N_1043),
	.LO(reg1_16[8])
);
defparam \d_cnst_sn.reg0_28_6_RNIKKH35_0[8] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNI6AH35_0[6]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg1_1 [6]),
	.I4(t_1[6]),
	.I5(N_1041),
	.LO(reg1_16[6])
);
defparam \d_cnst_sn.reg0_28_6_RNI6AH35_0[6] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNIR6095[5]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg0_1 [5]),
	.I4(t_1[5]),
	.I5(N_1040),
	.LO(reg0_28[5])
);
defparam \d_cnst_sn.reg0_28_6_RNIR6095[5] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNI6AH35[6]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg0_1 [6]),
	.I4(t_1[6]),
	.I5(N_1041),
	.LO(reg0_28[6])
);
defparam \d_cnst_sn.reg0_28_6_RNI6AH35[6] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNI9JV45[4]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg1_1 [4]),
	.I4(t_1[4]),
	.I5(N_1039),
	.LO(reg1_16[4])
);
defparam \d_cnst_sn.reg0_28_6_RNI9JV45[4] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNIR6095_0[5]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg1_1 [5]),
	.I4(t_1[5]),
	.I5(N_1040),
	.LO(reg1_16[5])
);
defparam \d_cnst_sn.reg0_28_6_RNIR6095_0[5] .INIT=64'h0F00FF0001001100;
// @7:74
  LUT6_L \d_cnst_sn.reg0_28_6_RNI9JV45_0[4]  (
	.I0(\d_cnst_sn.b64_0 ),
	.I1(\d_cnst_sn.b60_0 ),
	.I2(\d_cnst_sn.reg1_16_a0_1 [3]),
	.I3(\d_cnst_sn.reg0_1 [4]),
	.I4(t_1[4]),
	.I5(N_1039),
	.LO(reg0_28[4])
);
defparam \d_cnst_sn.reg0_28_6_RNI9JV45_0[4] .INIT=64'h0F00FF0001001100;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_5_RNIRBMC9[4]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_1_sqmuxa_RNIEMUH1),
	.I4(N_1816),
	.I5(r_4_2_a1_lut6_2_RNI2T8R3[3]),
	.LO(reg3_17[4])
);
defparam \d_cnst_sn.reg3_17_5_RNIRBMC9[4] .INIT=64'h777F0008F7FF8088;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_5_RNI2FMC9[5]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_1_sqmuxa_RNIHMUH1),
	.I4(N_1817),
	.I5(r_4_2_a1_lut6_2_RNI5V8R3[3]),
	.LO(reg3_17[5])
);
defparam \d_cnst_sn.reg3_17_5_RNI2FMC9[5] .INIT=64'h777F0008F7FF8088;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_5_RNIH8LK6[7]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_1_sqmuxa_RNINMUH1),
	.I4(N_1819),
	.I5(r_4_1_RNICM731[6]),
	.LO(reg3_17[7])
);
defparam \d_cnst_sn.reg3_17_5_RNIH8LK6[7] .INIT=64'h777F0008F7FF8088;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_5_RNIA5LK6[6]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_1_sqmuxa_RNIKMUH1),
	.I4(N_1818),
	.I5(r_4_1_RNI9K731[5]),
	.LO(reg3_17[6])
);
defparam \d_cnst_sn.reg3_17_5_RNIA5LK6[6] .INIT=64'h777F0008F7FF8088;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_5_RNIVELK6[9]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_1_sqmuxa_RNITMUH1),
	.I4(N_1821),
	.I5(r_4_1_RNIIQ731[8]),
	.LO(reg3_17[9])
);
defparam \d_cnst_sn.reg3_17_5_RNIVELK6[9] .INIT=64'h777F0008F7FF8088;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_5_RNIOBLK6[8]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_1_sqmuxa_RNIQMUH1),
	.I4(N_1820),
	.I5(r_4_1_RNIFO731[7]),
	.LO(reg3_17[8])
);
defparam \d_cnst_sn.reg3_17_5_RNIOBLK6[8] .INIT=64'h777F0008F7FF8088;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_5_RNI2DVL6[10]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_1_sqmuxa_RNIE1DM1),
	.I4(N_1822),
	.I5(r_4_1_RNIS3K91[9]),
	.LO(reg3_17[10])
);
defparam \d_cnst_sn.reg3_17_5_RNI2DVL6[10] .INIT=64'h777F0008F7FF8088;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_5_RNINL3U6[11]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_1_sqmuxa_RNIH1DM1),
	.I4(N_1823),
	.I5(r_4_1_RNIDBOH1[10]),
	.LO(reg3_17[11])
);
defparam \d_cnst_sn.reg3_17_5_RNINL3U6[11] .INIT=64'h777F0008F7FF8088;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[13]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(N_1670),
	.I3(\d_cnst_sn.reg3_17_6_1 [13]),
	.I4(N_1732),
	.I5(reg3_17_4_a2[13]),
	.LO(reg3_17[13])
);
defparam \d_cnst_sn.reg3_17[13] .INIT=64'h75752020FD75A820;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[27]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(\d_cnst_sn.reg3_17_6_0 [27]),
	.I3(N_1841),
	.I4(t_1[27]),
	.I5(N_1839),
	.LO(reg3_17[27])
);
defparam \d_cnst_sn.reg3_17[27] .INIT=64'hF0FFF4FFF000F400;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[28]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(\d_cnst_sn.reg3_17_6_0 [28]),
	.I3(N_1841),
	.I4(t_1[28]),
	.I5(N_1840),
	.LO(reg3_17[28])
);
defparam \d_cnst_sn.reg3_17[28] .INIT=64'hF0FFF4FFF000F400;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[16]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(N_1841),
	.I3(\d_cnst_sn.reg3_17_6_1 [16]),
	.I4(t_1[16]),
	.I5(N_1828),
	.LO(reg3_17[16])
);
defparam \d_cnst_sn.reg3_17[16] .INIT=64'hBF0FFF0FB000F000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[19]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(N_1841),
	.I3(\d_cnst_sn.reg3_17_6_1 [19]),
	.I4(t_1[19]),
	.I5(N_1831),
	.LO(reg3_17[19])
);
defparam \d_cnst_sn.reg3_17[19] .INIT=64'hBF0FFF0FB000F000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[20]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(\d_cnst_sn.reg3_17_6_0 [20]),
	.I3(N_1841),
	.I4(t_1[20]),
	.I5(N_1832),
	.LO(reg3_17[20])
);
defparam \d_cnst_sn.reg3_17[20] .INIT=64'hF0FFF4FFF000F400;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[14]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(t_1[14]),
	.I3(N_1841),
	.I4(\d_cnst_sn.reg3_17_6_1 [14]),
	.I5(N_1826),
	.LO(reg3_17[14])
);
defparam \d_cnst_sn.reg3_17[14] .INIT=64'hBFFF00FFBF000000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[18]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(N_1841),
	.I3(\d_cnst_sn.reg3_17_6_1 [18]),
	.I4(t_1[18]),
	.I5(N_1830),
	.LO(reg3_17[18])
);
defparam \d_cnst_sn.reg3_17[18] .INIT=64'hBF0FFF0FB000F000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[12]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(t_1[12]),
	.I3(N_1841),
	.I4(\d_cnst_sn.reg3_17_6_1 [12]),
	.I5(N_1824),
	.LO(reg3_17[12])
);
defparam \d_cnst_sn.reg3_17[12] .INIT=64'hBFFF00FFBF000000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[17]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(N_1841),
	.I3(\d_cnst_sn.reg3_17_6_1 [17]),
	.I4(t_1[17]),
	.I5(N_1829),
	.LO(reg3_17[17])
);
defparam \d_cnst_sn.reg3_17[17] .INIT=64'hBF0FFF0FB000F000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[15]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(N_1841),
	.I3(\d_cnst_sn.reg3_17_6_1 [15]),
	.I4(t_1[15]),
	.I5(N_1827),
	.LO(reg3_17[15])
);
defparam \d_cnst_sn.reg3_17[15] .INIT=64'hBF0FFF0FB000F000;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[26]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(\d_cnst_sn.reg3_17_6_0 [26]),
	.I3(N_1841),
	.I4(t_1[26]),
	.I5(N_1838),
	.LO(reg3_17[26])
);
defparam \d_cnst_sn.reg3_17[26] .INIT=64'hF0FFF4FFF000F400;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17[25]  (
	.I0(N_527_i),
	.I1(reg3_14_sqmuxa),
	.I2(\d_cnst_sn.reg3_17_6_0 [25]),
	.I3(N_1841),
	.I4(t_1[25]),
	.I5(N_1837),
	.LO(reg3_17[25])
);
defparam \d_cnst_sn.reg3_17[25] .INIT=64'hF0FFF4FFF000F400;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_2_RNI79973[24]  (
	.I0(N_1810),
	.I1(reg3_17_a0[24]),
	.I2(\d_cnst_sn.reg3_17_a1_2 [24]),
	.I3(\d_cnst_sn.reg3_17_0_tz [24]),
	.I4(t_1[24]),
	.I5(N_1743),
	.LO(reg3_17[24])
);
defparam \d_cnst_sn.reg3_17_2_RNI79973[24] .INIT=64'hFFDDFFFDEECCFEFC;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_2_RNI36973[23]  (
	.I0(N_1810),
	.I1(reg3_17_a0[23]),
	.I2(\d_cnst_sn.reg3_17_a1_2 [24]),
	.I3(\d_cnst_sn.reg3_17_0_tz [23]),
	.I4(t_1[23]),
	.I5(N_1742),
	.LO(reg3_17[23])
);
defparam \d_cnst_sn.reg3_17_2_RNI36973[23] .INIT=64'hFFDDFFFDEECCFEFC;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_2_RNIV2973[22]  (
	.I0(N_1810),
	.I1(reg3_17_a0[22]),
	.I2(\d_cnst_sn.reg3_17_a1_2 [24]),
	.I3(\d_cnst_sn.reg3_17_0_tz [22]),
	.I4(t_1[22]),
	.I5(N_1741),
	.LO(reg3_17[22])
);
defparam \d_cnst_sn.reg3_17_2_RNIV2973[22] .INIT=64'hFFDDFFFDEECCFEFC;
// @7:103
  LUT6_L \d_cnst_sn.reg3_17_2_RNIRV873[21]  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_0_tz [21]),
	.I2(reg3_17_a0[21]),
	.I3(\d_cnst_sn.reg3_17_a1_2 [24]),
	.I4(t_1[21]),
	.I5(N_1740),
	.LO(reg3_17[21])
);
defparam \d_cnst_sn.reg3_17_2_RNIRV873[21] .INIT=64'hFDFDFFFDF8F8FFF8;
// @7:47
  LUT6_L \d_cnst_sn.reg3_N_7_i_cZ  (
	.I0(N_1810),
	.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),
	.I2(reg3_14_sqmuxa),
	.I3(reg3_N_7_i_RNO),
	.I4(N_1815),
	.I5(t_6[3]),
	.LO(\d_cnst_sn.reg3_N_7_i )
);
defparam \d_cnst_sn.reg3_N_7_i_cZ .INIT=64'hF7FF8088777F0008;
  LUT5 \datai_RNI2IEL2[20]  (
	.I0(datai[20]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[20]),
	.O(un11_reg0_axb_20)
);
defparam \datai_RNI2IEL2[20] .INIT=32'hDDDF2220;
  LUT4 \datai_RNI2UAU_0[20]  (
	.I0(datai[20]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[20])
);
defparam \datai_RNI2UAU_0[20] .INIT=16'h2220;
  LUT5 \datai_RNIH7MC2[21]  (
	.I0(datai[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[21]),
	.O(un11_reg0_axb_21)
);
defparam \datai_RNIH7MC2[21] .INIT=32'hDDDF2220;
  LUT4 \datai_RNI3VAU_0[21]  (
	.I0(datai[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[21])
);
defparam \datai_RNI3VAU_0[21] .INIT=16'h2220;
  LUT5 \datai_RNIAOEL2[22]  (
	.I0(datai[22]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[22]),
	.O(un11_reg0_axb_22)
);
defparam \datai_RNIAOEL2[22] .INIT=32'hDDDF2220;
  LUT4 \datai_RNI40BU_0[22]  (
	.I0(datai[22]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[22])
);
defparam \datai_RNI40BU_0[22] .INIT=16'h2220;
  LUT5 \datai_RNI5SEL2[23]  (
	.I0(datai[23]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[23]),
	.O(un11_reg0_axb_23)
);
defparam \datai_RNI5SEL2[23] .INIT=32'hDDDF2220;
  LUT4 \datai_RNI51BU_0[23]  (
	.I0(datai[23]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[23])
);
defparam \datai_RNI51BU_0[23] .INIT=16'h2220;
  LUT5 \datai_RNI9VEL2[24]  (
	.I0(datai[24]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[24]),
	.O(un11_reg0_axb_24)
);
defparam \datai_RNI9VEL2[24] .INIT=32'hDDDF2220;
  LUT4 \datai_RNI62BU_0[24]  (
	.I0(datai[24]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[24])
);
defparam \datai_RNI62BU_0[24] .INIT=16'h2220;
  LUT5 \datai_RNI1OMC2[25]  (
	.I0(datai[25]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[25]),
	.O(un11_reg0_axb_25)
);
defparam \datai_RNI1OMC2[25] .INIT=32'hDDDF2220;
  LUT4 \datai_RNI73BU_0[25]  (
	.I0(datai[25]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[25])
);
defparam \datai_RNI73BU_0[25] .INIT=16'h2220;
  LUT5 \datai_RNI5SMC2[26]  (
	.I0(datai[26]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[26]),
	.O(un11_reg0_axb_26)
);
defparam \datai_RNI5SMC2[26] .INIT=32'hDDDF2220;
  LUT4 \datai_RNI84BU_0[26]  (
	.I0(datai[26]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[26])
);
defparam \datai_RNI84BU_0[26] .INIT=16'h2220;
  LUT5 \datai_RNIL8FL2[27]  (
	.I0(datai[27]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[27]),
	.O(un11_reg0_axb_27)
);
defparam \datai_RNIL8FL2[27] .INIT=32'hDDDF2220;
  LUT4 \datai_RNI95BU_0[27]  (
	.I0(datai[27]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[27])
);
defparam \datai_RNI95BU_0[27] .INIT=16'h2220;
  LUT5 \datai_RNID4NC2[28]  (
	.I0(datai[28]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.I4(r_4[28]),
	.O(un11_reg0_axb_28)
);
defparam \datai_RNID4NC2[28] .INIT=32'hDDDF2220;
  LUT4 \datai_RNIA6BU_0[28]  (
	.I0(datai[28]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[28])
);
defparam \datai_RNIA6BU_0[28] .INIT=16'h2220;
  LUT5 \d_cnst_sn.r_4_1_RNI4OE61[5]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_920),
	.I3(N_952),
	.I4(m_2[5]),
	.O(un32_reg0_axb_5)
);
defparam \d_cnst_sn.r_4_1_RNI4OE61[5] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNI7RE61[6]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_921),
	.I3(N_953),
	.I4(m_2[6]),
	.O(un32_reg0_axb_6)
);
defparam \d_cnst_sn.r_4_1_RNI7RE61[6] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNIAUE61[7]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_922),
	.I3(N_954),
	.I4(m_2[7]),
	.O(un32_reg0_axb_7)
);
defparam \d_cnst_sn.r_4_1_RNIAUE61[7] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNID1F61[8]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_923),
	.I3(N_955),
	.I4(m_2[8]),
	.O(un32_reg0_axb_8)
);
defparam \d_cnst_sn.r_4_1_RNID1F61[8] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNIG4F61[9]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_924),
	.I3(N_956),
	.I4(m_2[9]),
	.O(un32_reg0_axb_9)
);
defparam \d_cnst_sn.r_4_1_RNIG4F61[9] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNI88L31[10]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_925),
	.I3(N_957),
	.I4(m_2[10]),
	.O(un32_reg0_axb_10)
);
defparam \d_cnst_sn.r_4_1_RNI88L31[10] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNIBBL31[11]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_926),
	.I3(N_958),
	.I4(m_2[11]),
	.O(un32_reg0_axb_11)
);
defparam \d_cnst_sn.r_4_1_RNIBBL31[11] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNIEEL31[12]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_927),
	.I3(N_959),
	.I4(m_2[12]),
	.O(un32_reg0_axb_12)
);
defparam \d_cnst_sn.r_4_1_RNIEEL31[12] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNIHHL31[13]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_928),
	.I3(N_960),
	.I4(m_2[13]),
	.O(un32_reg0_axb_13)
);
defparam \d_cnst_sn.r_4_1_RNIHHL31[13] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNIKKL31[14]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_929),
	.I3(N_961),
	.I4(m_2[14]),
	.O(un32_reg0_axb_14)
);
defparam \d_cnst_sn.r_4_1_RNIKKL31[14] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNINNL31[15]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_930),
	.I3(N_962),
	.I4(m_2[15]),
	.O(un32_reg0_axb_15)
);
defparam \d_cnst_sn.r_4_1_RNINNL31[15] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNIQQL31[16]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_931),
	.I3(N_963),
	.I4(m_2[16]),
	.O(un32_reg0_axb_16)
);
defparam \d_cnst_sn.r_4_1_RNIQQL31[16] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNITTL31[17]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_932),
	.I3(N_964),
	.I4(m_2[17]),
	.O(un32_reg0_axb_17)
);
defparam \d_cnst_sn.r_4_1_RNITTL31[17] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNI01M31[18]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_933),
	.I3(N_965),
	.I4(m_2[18]),
	.O(un32_reg0_axb_18)
);
defparam \d_cnst_sn.r_4_1_RNI01M31[18] .INIT=32'hF4B00B4F;
  LUT5 \d_cnst_sn.r_4_1_RNIOJPQ1[19]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[29]),
	.I2(N_934),
	.I3(N_2722),
	.I4(m_2[19]),
	.O(un32_reg0_axb_19)
);
defparam \d_cnst_sn.r_4_1_RNIOJPQ1[19] .INIT=32'hF4B00B4F;
// @7:466
  XORCY t_1_s_31 (
	.LI(r_4[31]),
	.CI(t_1_cry_30),
	.O(t_1[31])
);
// @7:466
  XORCY t_1_s_30 (
	.LI(N_4571_i),
	.CI(t_1_cry_29),
	.O(t_1[30])
);
// @7:466
  MUXCY_L t_1_cry_30_cZ (
	.DI(VCC),
	.CI(t_1_cry_29),
	.S(N_4571_i),
	.LO(t_1_cry_30)
);
// @7:466
  XORCY t_1_s_29 (
	.LI(N_4570_i),
	.CI(t_1_cry_28),
	.O(t_1[29])
);
// @7:466
  MUXCY_L t_1_cry_29_cZ (
	.DI(VCC),
	.CI(t_1_cry_28),
	.S(N_4570_i),
	.LO(t_1_cry_29)
);
// @7:466
  XORCY t_1_s_28 (
	.LI(N_4569_i),
	.CI(t_1_cry_27),
	.O(t_1[28])
);
// @7:466
  MUXCY_L t_1_cry_28_cZ (
	.DI(VCC),
	.CI(t_1_cry_27),
	.S(N_4569_i),
	.LO(t_1_cry_28)
);
// @7:466
  XORCY t_1_s_27 (
	.LI(N_4568_i),
	.CI(t_1_cry_26),
	.O(t_1[27])
);
// @7:466
  MUXCY_L t_1_cry_27_cZ (
	.DI(VCC),
	.CI(t_1_cry_26),
	.S(N_4568_i),
	.LO(t_1_cry_27)
);
// @7:466
  XORCY t_1_s_26 (
	.LI(N_4567_i),
	.CI(t_1_cry_25),
	.O(t_1[26])
);
// @7:466
  MUXCY_L t_1_cry_26_cZ (
	.DI(VCC),
	.CI(t_1_cry_25),
	.S(N_4567_i),
	.LO(t_1_cry_26)
);
// @7:466
  XORCY t_1_s_25 (
	.LI(N_4566_i),
	.CI(t_1_cry_24),
	.O(t_1[25])
);
// @7:466
  MUXCY_L t_1_cry_25_cZ (
	.DI(VCC),
	.CI(t_1_cry_24),
	.S(N_4566_i),
	.LO(t_1_cry_25)
);
// @7:466
  XORCY t_1_s_24 (
	.LI(N_4565_i),
	.CI(t_1_cry_23),
	.O(t_1[24])
);
// @7:466
  MUXCY_L t_1_cry_24_cZ (
	.DI(VCC),
	.CI(t_1_cry_23),
	.S(N_4565_i),
	.LO(t_1_cry_24)
);
// @7:466
  XORCY t_1_s_23 (
	.LI(N_4564_i),
	.CI(t_1_cry_22),
	.O(t_1[23])
);
// @7:466
  MUXCY_L t_1_cry_23_cZ (
	.DI(VCC),
	.CI(t_1_cry_22),
	.S(N_4564_i),
	.LO(t_1_cry_23)
);
// @7:466
  XORCY t_1_s_22 (
	.LI(N_4563_i),
	.CI(t_1_cry_21),
	.O(t_1[22])
);
// @7:466
  MUXCY_L t_1_cry_22_cZ (
	.DI(VCC),
	.CI(t_1_cry_21),
	.S(N_4563_i),
	.LO(t_1_cry_22)
);
// @7:466
  XORCY t_1_s_21 (
	.LI(N_4562_i),
	.CI(t_1_cry_20),
	.O(t_1[21])
);
// @7:466
  MUXCY_L t_1_cry_21_cZ (
	.DI(VCC),
	.CI(t_1_cry_20),
	.S(N_4562_i),
	.LO(t_1_cry_21)
);
// @7:466
  XORCY t_1_s_20 (
	.LI(N_4561_i),
	.CI(t_1_cry_19),
	.O(t_1[20])
);
// @7:466
  MUXCY_L t_1_cry_20_cZ (
	.DI(VCC),
	.CI(t_1_cry_19),
	.S(N_4561_i),
	.LO(t_1_cry_20)
);
// @7:466
  XORCY t_1_s_19 (
	.LI(N_4560_i),
	.CI(t_1_cry_18),
	.O(t_1[19])
);
// @7:466
  MUXCY_L t_1_cry_19_cZ (
	.DI(VCC),
	.CI(t_1_cry_18),
	.S(N_4560_i),
	.LO(t_1_cry_19)
);
// @7:466
  XORCY t_1_s_18 (
	.LI(N_4559_i),
	.CI(t_1_cry_17),
	.O(t_1[18])
);
// @7:466
  MUXCY_L t_1_cry_18_cZ (
	.DI(VCC),
	.CI(t_1_cry_17),
	.S(N_4559_i),
	.LO(t_1_cry_18)
);
// @7:466
  XORCY t_1_s_17 (
	.LI(N_4558_i),
	.CI(t_1_cry_16),
	.O(t_1[17])
);
// @7:466
  MUXCY_L t_1_cry_17_cZ (
	.DI(VCC),
	.CI(t_1_cry_16),
	.S(N_4558_i),
	.LO(t_1_cry_17)
);
// @7:466
  XORCY t_1_s_16 (
	.LI(N_4557_i),
	.CI(t_1_cry_15),
	.O(t_1[16])
);
// @7:466
  MUXCY_L t_1_cry_16_cZ (
	.DI(VCC),
	.CI(t_1_cry_15),
	.S(N_4557_i),
	.LO(t_1_cry_16)
);
// @7:466
  XORCY t_1_s_15 (
	.LI(N_4556_i),
	.CI(t_1_cry_14),
	.O(t_1[15])
);
// @7:466
  MUXCY_L t_1_cry_15_cZ (
	.DI(VCC),
	.CI(t_1_cry_14),
	.S(N_4556_i),
	.LO(t_1_cry_15)
);
// @7:466
  XORCY t_1_s_14 (
	.LI(N_4555_i),
	.CI(t_1_cry_13),
	.O(t_1[14])
);
// @7:466
  MUXCY_L t_1_cry_14_cZ (
	.DI(VCC),
	.CI(t_1_cry_13),
	.S(N_4555_i),
	.LO(t_1_cry_14)
);
// @7:466
  XORCY t_1_s_13 (
	.LI(N_4554_i),
	.CI(t_1_cry_12),
	.O(t_1[13])
);
// @7:466
  MUXCY_L t_1_cry_13_cZ (
	.DI(VCC),
	.CI(t_1_cry_12),
	.S(N_4554_i),
	.LO(t_1_cry_13)
);
// @7:466
  XORCY t_1_s_12 (
	.LI(N_4553_i),
	.CI(t_1_cry_11),
	.O(t_1[12])
);
// @7:466
  MUXCY_L t_1_cry_12_cZ (
	.DI(VCC),
	.CI(t_1_cry_11),
	.S(N_4553_i),
	.LO(t_1_cry_12)
);
// @7:466
  XORCY t_1_s_11 (
	.LI(N_4552_i),
	.CI(t_1_cry_10),
	.O(t_1[11])
);
// @7:466
  MUXCY_L t_1_cry_11_cZ (
	.DI(VCC),
	.CI(t_1_cry_10),
	.S(N_4552_i),
	.LO(t_1_cry_11)
);
// @7:466
  XORCY t_1_s_10 (
	.LI(N_4551_i),
	.CI(t_1_cry_9),
	.O(t_1[10])
);
// @7:466
  MUXCY_L t_1_cry_10_cZ (
	.DI(VCC),
	.CI(t_1_cry_9),
	.S(N_4551_i),
	.LO(t_1_cry_10)
);
// @7:466
  XORCY t_1_s_9 (
	.LI(N_4550_i),
	.CI(t_1_cry_8),
	.O(t_1[9])
);
// @7:466
  MUXCY_L t_1_cry_9_cZ (
	.DI(VCC),
	.CI(t_1_cry_8),
	.S(N_4550_i),
	.LO(t_1_cry_9)
);
// @7:466
  XORCY t_1_s_8 (
	.LI(N_4549_i),
	.CI(t_1_cry_7),
	.O(t_1[8])
);
// @7:466
  MUXCY_L t_1_cry_8_cZ (
	.DI(VCC),
	.CI(t_1_cry_7),
	.S(N_4549_i),
	.LO(t_1_cry_8)
);
// @7:466
  XORCY t_1_s_7 (
	.LI(N_4548_i),
	.CI(t_1_cry_6),
	.O(t_1[7])
);
// @7:466
  MUXCY_L t_1_cry_7_cZ (
	.DI(VCC),
	.CI(t_1_cry_6),
	.S(N_4548_i),
	.LO(t_1_cry_7)
);
// @7:466
  XORCY t_1_s_6 (
	.LI(N_4547_i),
	.CI(t_1_cry_5),
	.O(t_1[6])
);
// @7:466
  MUXCY_L t_1_cry_6_cZ (
	.DI(VCC),
	.CI(t_1_cry_5),
	.S(N_4547_i),
	.LO(t_1_cry_6)
);
// @7:466
  XORCY t_1_s_5 (
	.LI(N_4546_i),
	.CI(t_1_cry_4),
	.O(t_1[5])
);
// @7:466
  MUXCY_L t_1_cry_5_cZ (
	.DI(VCC),
	.CI(t_1_cry_4),
	.S(N_4546_i),
	.LO(t_1_cry_5)
);
// @7:466
  XORCY t_1_s_4 (
	.LI(N_4545_i),
	.CI(t_1_cry_3),
	.O(t_1[4])
);
// @7:466
  MUXCY_L t_1_cry_4_cZ (
	.DI(VCC),
	.CI(t_1_cry_3),
	.S(N_4545_i),
	.LO(t_1_cry_4)
);
// @7:466
  XORCY t_1_s_3 (
	.LI(N_4544_i),
	.CI(t_1_cry_2),
	.O(t_1[3])
);
// @7:466
  MUXCY_L t_1_cry_3_cZ (
	.DI(VCC),
	.CI(t_1_cry_2),
	.S(N_4544_i),
	.LO(t_1_cry_3)
);
// @7:466
  XORCY t_1_s_2 (
	.LI(N_4543_i),
	.CI(t_1_cry_1),
	.O(t_1[2])
);
// @7:466
  MUXCY_L t_1_cry_2_cZ (
	.DI(VCC),
	.CI(t_1_cry_1),
	.S(N_4543_i),
	.LO(t_1_cry_2)
);
// @7:466
  XORCY t_1_s_1 (
	.LI(N_4542_i),
	.CI(t_1_cry_0),
	.O(t_1[1])
);
// @7:466
  MUXCY_L t_1_cry_1_cZ (
	.DI(VCC),
	.CI(t_1_cry_0),
	.S(N_4542_i),
	.LO(t_1_cry_1)
);
// @7:466
  XORCY t_1_s_0 (
	.LI(N_4541_i),
	.CI(t_1_cry_0_cy),
	.O(t_1[0])
);
// @7:466
  MUXCY_L t_1_cry_0_cZ (
	.DI(VCC),
	.CI(t_1_cry_0_cy),
	.S(N_4541_i),
	.LO(t_1_cry_0)
);
// @7:95
  XORCY un3_reg3_s_25_cZ (
	.LI(un3_reg3_axb_25),
	.CI(un3_reg3_cry_24),
	.O(un3_reg3_s_25)
);
// @7:95
  MUXCY un3_reg3_cry_25_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_24),
	.S(un3_reg3_axb_25),
	.O(un3_reg3_cry_25_0)
);
// @7:95
  XORCY un3_reg3_s_24_cZ (
	.LI(un3_reg3_axb_24),
	.CI(un3_reg3_cry_23),
	.O(un3_reg3_s_24)
);
// @7:95
  MUXCY_L un3_reg3_cry_24_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_23),
	.S(un3_reg3_axb_24),
	.LO(un3_reg3_cry_24)
);
// @7:95
  XORCY un3_reg3_s_23_cZ (
	.LI(un3_reg3_axb_23),
	.CI(un3_reg3_cry_22),
	.O(un3_reg3_s_23)
);
// @7:95
  MUXCY_L un3_reg3_cry_23_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_22),
	.S(un3_reg3_axb_23),
	.LO(un3_reg3_cry_23)
);
// @7:95
  XORCY un3_reg3_s_22_cZ (
	.LI(un3_reg3_axb_22),
	.CI(un3_reg3_cry_21),
	.O(un3_reg3_s_22)
);
// @7:95
  MUXCY_L un3_reg3_cry_22_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_21),
	.S(un3_reg3_axb_22),
	.LO(un3_reg3_cry_22)
);
// @7:95
  XORCY un3_reg3_s_21_cZ (
	.LI(un3_reg3_axb_21),
	.CI(un3_reg3_cry_20),
	.O(un3_reg3_s_21)
);
// @7:95
  MUXCY_L un3_reg3_cry_21_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_20),
	.S(un3_reg3_axb_21),
	.LO(un3_reg3_cry_21)
);
// @7:95
  XORCY un3_reg3_s_20_cZ (
	.LI(un3_reg3_axb_20),
	.CI(un3_reg3_cry_19),
	.O(un3_reg3_s_20)
);
// @7:95
  MUXCY_L un3_reg3_cry_20_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_19),
	.S(un3_reg3_axb_20),
	.LO(un3_reg3_cry_20)
);
// @7:95
  XORCY un3_reg3_s_19_cZ (
	.LI(un3_reg3_axb_19),
	.CI(un3_reg3_cry_18),
	.O(un3_reg3_s_19)
);
// @7:95
  MUXCY_L un3_reg3_cry_19_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_18),
	.S(un3_reg3_axb_19),
	.LO(un3_reg3_cry_19)
);
// @7:95
  XORCY un3_reg3_s_18_cZ (
	.LI(un3_reg3_axb_18),
	.CI(un3_reg3_cry_17),
	.O(un3_reg3_s_18)
);
// @7:95
  MUXCY_L un3_reg3_cry_18_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_17),
	.S(un3_reg3_axb_18),
	.LO(un3_reg3_cry_18)
);
// @7:95
  XORCY un3_reg3_s_17_cZ (
	.LI(un3_reg3_axb_17),
	.CI(un3_reg3_cry_16),
	.O(un3_reg3_s_17)
);
// @7:95
  MUXCY_L un3_reg3_cry_17_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_16),
	.S(un3_reg3_axb_17),
	.LO(un3_reg3_cry_17)
);
// @7:95
  XORCY un3_reg3_s_16_cZ (
	.LI(un3_reg3_axb_16),
	.CI(un3_reg3_cry_15),
	.O(un3_reg3_s_16)
);
// @7:95
  MUXCY_L un3_reg3_cry_16_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_15),
	.S(un3_reg3_axb_16),
	.LO(un3_reg3_cry_16)
);
// @7:95
  XORCY un3_reg3_s_15_cZ (
	.LI(un3_reg3_axb_15),
	.CI(un3_reg3_cry_14),
	.O(un3_reg3_s_15)
);
// @7:95
  MUXCY_L un3_reg3_cry_15_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_14),
	.S(un3_reg3_axb_15),
	.LO(un3_reg3_cry_15)
);
// @7:95
  XORCY un3_reg3_s_14_cZ (
	.LI(un3_reg3_axb_14),
	.CI(un3_reg3_cry_13),
	.O(un3_reg3_s_14)
);
// @7:95
  MUXCY_L un3_reg3_cry_14_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_13),
	.S(un3_reg3_axb_14),
	.LO(un3_reg3_cry_14)
);
// @7:95
  XORCY un3_reg3_s_13_cZ (
	.LI(un3_reg3_axb_13),
	.CI(un3_reg3_cry_12),
	.O(un3_reg3_s_13)
);
// @7:95
  MUXCY_L un3_reg3_cry_13_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_12),
	.S(un3_reg3_axb_13),
	.LO(un3_reg3_cry_13)
);
// @7:95
  XORCY un3_reg3_s_12_cZ (
	.LI(un3_reg3_axb_12),
	.CI(un3_reg3_cry_11),
	.O(un3_reg3_s_12)
);
// @7:95
  MUXCY_L un3_reg3_cry_12_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_11),
	.S(un3_reg3_axb_12),
	.LO(un3_reg3_cry_12)
);
// @7:95
  XORCY un3_reg3_s_11_cZ (
	.LI(un3_reg3_axb_11),
	.CI(un3_reg3_cry_10),
	.O(un3_reg3_s_11)
);
// @7:95
  MUXCY_L un3_reg3_cry_11_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_10),
	.S(un3_reg3_axb_11),
	.LO(un3_reg3_cry_11)
);
// @7:95
  XORCY un3_reg3_s_10_cZ (
	.LI(un3_reg3_axb_10),
	.CI(un3_reg3_cry_9),
	.O(un3_reg3_s_10)
);
// @7:95
  MUXCY_L un3_reg3_cry_10_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_9),
	.S(un3_reg3_axb_10),
	.LO(un3_reg3_cry_10)
);
// @7:95
  XORCY un3_reg3_s_9_cZ (
	.LI(un3_reg3_axb_9),
	.CI(un3_reg3_cry_8),
	.O(un3_reg3_s_9)
);
// @7:95
  MUXCY_L un3_reg3_cry_9_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_8),
	.S(un3_reg3_axb_9),
	.LO(un3_reg3_cry_9)
);
// @7:95
  XORCY un3_reg3_s_8_cZ (
	.LI(un3_reg3_axb_8),
	.CI(un3_reg3_cry_7),
	.O(un3_reg3_s_8)
);
// @7:95
  MUXCY_L un3_reg3_cry_8_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_7),
	.S(un3_reg3_axb_8),
	.LO(un3_reg3_cry_8)
);
// @7:95
  XORCY un3_reg3_s_7_cZ (
	.LI(un3_reg3_axb_7),
	.CI(un3_reg3_cry_6),
	.O(un3_reg3_s_7)
);
// @7:95
  MUXCY_L un3_reg3_cry_7_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_6),
	.S(un3_reg3_axb_7),
	.LO(un3_reg3_cry_7)
);
// @7:95
  XORCY un3_reg3_s_6_cZ (
	.LI(un3_reg3_axb_6),
	.CI(un3_reg3_cry_5),
	.O(un3_reg3_s_6)
);
// @7:95
  MUXCY_L un3_reg3_cry_6_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_5),
	.S(un3_reg3_axb_6),
	.LO(un3_reg3_cry_6)
);
// @7:95
  XORCY un3_reg3_s_5_cZ (
	.LI(un3_reg3_axb_5),
	.CI(un3_reg3_cry_4),
	.O(un3_reg3_s_5)
);
// @7:95
  MUXCY_L un3_reg3_cry_5_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_4),
	.S(un3_reg3_axb_5),
	.LO(un3_reg3_cry_5)
);
// @7:95
  XORCY un3_reg3_s_4_cZ (
	.LI(un3_reg3_axb_4),
	.CI(un3_reg3_cry_3),
	.O(un3_reg3_s_4)
);
// @7:95
  MUXCY_L un3_reg3_cry_4_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_3),
	.S(un3_reg3_axb_4),
	.LO(un3_reg3_cry_4)
);
// @7:95
  XORCY un3_reg3_s_3_cZ (
	.LI(un3_reg3_axb_3),
	.CI(un3_reg3_cry_2),
	.O(un3_reg3_s_3)
);
// @7:95
  MUXCY_L un3_reg3_cry_3_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_2),
	.S(un3_reg3_axb_3),
	.LO(un3_reg3_cry_3)
);
// @7:95
  XORCY un3_reg3_s_2_cZ (
	.LI(un3_reg3_axb_2),
	.CI(un3_reg3_cry_1),
	.O(un3_reg3_s_2)
);
// @7:95
  MUXCY_L un3_reg3_cry_2_cZ (
	.DI(GND),
	.CI(un3_reg3_cry_1),
	.S(un3_reg3_axb_2),
	.LO(un3_reg3_cry_2)
);
// @7:95
  XORCY un3_reg3_s_1_cZ (
	.LI(un3_reg3_axb_1),
	.CI(reg3[3]),
	.O(un3_reg3_s_1)
);
// @7:95
  MUXCY_L un3_reg3_cry_1_cZ (
	.DI(GND),
	.CI(reg3[3]),
	.S(un3_reg3_axb_1),
	.LO(un3_reg3_cry_1)
);
// @7:74
  XORCY un1_inf_abs0_0_s_19 (
	.LI(un1_inf_abs0_0_axb_19),
	.CI(un1_inf_abs0_0_cry_18),
	.O(un1_inf_abs0_11[19])
);
// @7:74
  XORCY un1_inf_abs0_0_s_18 (
	.LI(un1_inf_abs0_0_axb_18),
	.CI(un1_inf_abs0_0_cry_17),
	.O(un1_inf_abs0_11[18])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_18_cZ (
	.DI(inf_abs0_2[18]),
	.CI(un1_inf_abs0_0_cry_17),
	.S(un1_inf_abs0_0_axb_18),
	.LO(un1_inf_abs0_0_cry_18)
);
// @7:74
  XORCY un1_inf_abs0_0_s_17 (
	.LI(un1_inf_abs0_0_axb_17),
	.CI(un1_inf_abs0_0_cry_16),
	.O(un1_inf_abs0_11[17])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_17_cZ (
	.DI(inf_abs0_2[17]),
	.CI(un1_inf_abs0_0_cry_16),
	.S(un1_inf_abs0_0_axb_17),
	.LO(un1_inf_abs0_0_cry_17)
);
// @7:74
  XORCY un1_inf_abs0_0_s_16 (
	.LI(un1_inf_abs0_0_axb_16),
	.CI(un1_inf_abs0_0_cry_15),
	.O(un1_inf_abs0_11[16])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_16_cZ (
	.DI(inf_abs0_2[16]),
	.CI(un1_inf_abs0_0_cry_15),
	.S(un1_inf_abs0_0_axb_16),
	.LO(un1_inf_abs0_0_cry_16)
);
// @7:74
  XORCY un1_inf_abs0_0_s_15 (
	.LI(un1_inf_abs0_0_axb_15),
	.CI(un1_inf_abs0_0_cry_14),
	.O(un1_inf_abs0_11[15])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_15_cZ (
	.DI(inf_abs0_2[15]),
	.CI(un1_inf_abs0_0_cry_14),
	.S(un1_inf_abs0_0_axb_15),
	.LO(un1_inf_abs0_0_cry_15)
);
// @7:74
  XORCY un1_inf_abs0_0_s_14 (
	.LI(un1_inf_abs0_0_axb_14),
	.CI(un1_inf_abs0_0_cry_13),
	.O(un1_inf_abs0_11[14])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_14_cZ (
	.DI(inf_abs0_2[14]),
	.CI(un1_inf_abs0_0_cry_13),
	.S(un1_inf_abs0_0_axb_14),
	.LO(un1_inf_abs0_0_cry_14)
);
// @7:74
  XORCY un1_inf_abs0_0_s_13 (
	.LI(un1_inf_abs0_0_axb_13),
	.CI(un1_inf_abs0_0_cry_12),
	.O(un1_inf_abs0_11[13])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_13_cZ (
	.DI(inf_abs0_2[13]),
	.CI(un1_inf_abs0_0_cry_12),
	.S(un1_inf_abs0_0_axb_13),
	.LO(un1_inf_abs0_0_cry_13)
);
// @7:74
  XORCY un1_inf_abs0_0_s_12 (
	.LI(un1_inf_abs0_0_axb_12),
	.CI(un1_inf_abs0_0_cry_11),
	.O(un1_inf_abs0_11[12])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_12_cZ (
	.DI(inf_abs0_2[12]),
	.CI(un1_inf_abs0_0_cry_11),
	.S(un1_inf_abs0_0_axb_12),
	.LO(un1_inf_abs0_0_cry_12)
);
// @7:74
  XORCY un1_inf_abs0_0_s_11 (
	.LI(un1_inf_abs0_0_axb_11),
	.CI(un1_inf_abs0_0_cry_10),
	.O(un1_inf_abs0_11[11])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_11_cZ (
	.DI(inf_abs0_2[11]),
	.CI(un1_inf_abs0_0_cry_10),
	.S(un1_inf_abs0_0_axb_11),
	.LO(un1_inf_abs0_0_cry_11)
);
// @7:74
  XORCY un1_inf_abs0_0_s_10 (
	.LI(un1_inf_abs0_0_axb_10),
	.CI(un1_inf_abs0_0_cry_9),
	.O(un1_inf_abs0_11[10])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_10_cZ (
	.DI(inf_abs0_2[10]),
	.CI(un1_inf_abs0_0_cry_9),
	.S(un1_inf_abs0_0_axb_10),
	.LO(un1_inf_abs0_0_cry_10)
);
// @7:74
  XORCY un1_inf_abs0_0_s_9 (
	.LI(un1_inf_abs0_0_axb_9),
	.CI(un1_inf_abs0_0_cry_8),
	.O(un1_inf_abs0_11[9])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_9_cZ (
	.DI(inf_abs0_2[9]),
	.CI(un1_inf_abs0_0_cry_8),
	.S(un1_inf_abs0_0_axb_9),
	.LO(un1_inf_abs0_0_cry_9)
);
// @7:74
  XORCY un1_inf_abs0_0_s_8 (
	.LI(un1_inf_abs0_0_axb_8),
	.CI(un1_inf_abs0_0_cry_7),
	.O(un1_inf_abs0_11[8])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_8_cZ (
	.DI(inf_abs0_2[8]),
	.CI(un1_inf_abs0_0_cry_7),
	.S(un1_inf_abs0_0_axb_8),
	.LO(un1_inf_abs0_0_cry_8)
);
// @7:74
  XORCY un1_inf_abs0_0_s_7 (
	.LI(un1_inf_abs0_0_axb_7),
	.CI(un1_inf_abs0_0_cry_6),
	.O(un1_inf_abs0_11[7])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_7_cZ (
	.DI(inf_abs0_2[7]),
	.CI(un1_inf_abs0_0_cry_6),
	.S(un1_inf_abs0_0_axb_7),
	.LO(un1_inf_abs0_0_cry_7)
);
// @7:74
  XORCY un1_inf_abs0_0_s_6 (
	.LI(un1_inf_abs0_0_axb_6),
	.CI(un1_inf_abs0_0_cry_5),
	.O(un1_inf_abs0_11[6])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_6_cZ (
	.DI(inf_abs0_2[6]),
	.CI(un1_inf_abs0_0_cry_5),
	.S(un1_inf_abs0_0_axb_6),
	.LO(un1_inf_abs0_0_cry_6)
);
// @7:74
  XORCY un1_inf_abs0_0_s_5 (
	.LI(un1_inf_abs0_0_axb_5),
	.CI(un1_inf_abs0_0_cry_4),
	.O(un1_inf_abs0_11[5])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_5_cZ (
	.DI(inf_abs0_2[5]),
	.CI(un1_inf_abs0_0_cry_4),
	.S(un1_inf_abs0_0_axb_5),
	.LO(un1_inf_abs0_0_cry_5)
);
// @7:74
  XORCY un1_inf_abs0_0_s_4 (
	.LI(un1_inf_abs0_0_axb_4),
	.CI(un1_inf_abs0_0_cry_3),
	.O(un1_inf_abs0_11[4])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_4_cZ (
	.DI(inf_abs0_2[4]),
	.CI(un1_inf_abs0_0_cry_3),
	.S(un1_inf_abs0_0_axb_4),
	.LO(un1_inf_abs0_0_cry_4)
);
// @7:74
  XORCY un1_inf_abs0_0_s_3 (
	.LI(un1_inf_abs0_0_axb_3),
	.CI(un1_inf_abs0_0_cry_2),
	.O(un1_inf_abs0_11[3])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_3_cZ (
	.DI(inf_abs0_2[3]),
	.CI(un1_inf_abs0_0_cry_2),
	.S(un1_inf_abs0_0_axb_3),
	.LO(un1_inf_abs0_0_cry_3)
);
// @7:74
  XORCY un1_inf_abs0_0_s_2 (
	.LI(un1_inf_abs0_0_axb_2),
	.CI(un1_inf_abs0_0_cry_1),
	.O(un1_inf_abs0_11[2])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_2_cZ (
	.DI(inf_abs0_2[2]),
	.CI(un1_inf_abs0_0_cry_1),
	.S(un1_inf_abs0_0_axb_2),
	.LO(un1_inf_abs0_0_cry_2)
);
// @7:74
  XORCY un1_inf_abs0_0_s_1 (
	.LI(un1_inf_abs0_0_axb_1),
	.CI(un1_inf_abs0_0_cry_0),
	.O(un1_inf_abs0_11[1])
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_1_cZ (
	.DI(inf_abs0_2[1]),
	.CI(un1_inf_abs0_0_cry_0),
	.S(un1_inf_abs0_0_axb_1),
	.LO(un1_inf_abs0_0_cry_1)
);
// @7:74
  MUXCY_L un1_inf_abs0_0_cry_0_cZ (
	.DI(inf_abs0_2[0]),
	.CI(GND),
	.S(un1_inf_abs0_11[0]),
	.LO(un1_inf_abs0_0_cry_0)
);
// @7:74
  XORCY un1_inf_abs0_s_19 (
	.LI(un1_inf_abs0_axb_19),
	.CI(un1_inf_abs0_cry_18),
	.O(un1_inf_abs0_10[19])
);
// @7:74
  XORCY un1_inf_abs0_s_18 (
	.LI(un1_inf_abs0_axb_18),
	.CI(un1_inf_abs0_cry_17),
	.O(un1_inf_abs0_10[18])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_18_cZ (
	.DI(inf_abs0_2[18]),
	.CI(un1_inf_abs0_cry_17),
	.S(un1_inf_abs0_axb_18),
	.LO(un1_inf_abs0_cry_18)
);
// @7:74
  XORCY un1_inf_abs0_s_17 (
	.LI(un1_inf_abs0_axb_17),
	.CI(un1_inf_abs0_cry_16),
	.O(un1_inf_abs0_10[17])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_17_cZ (
	.DI(inf_abs0_2[17]),
	.CI(un1_inf_abs0_cry_16),
	.S(un1_inf_abs0_axb_17),
	.LO(un1_inf_abs0_cry_17)
);
// @7:74
  XORCY un1_inf_abs0_s_16 (
	.LI(un1_inf_abs0_axb_16),
	.CI(un1_inf_abs0_cry_15),
	.O(un1_inf_abs0_10[16])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_16_cZ (
	.DI(inf_abs0_2[16]),
	.CI(un1_inf_abs0_cry_15),
	.S(un1_inf_abs0_axb_16),
	.LO(un1_inf_abs0_cry_16)
);
// @7:74
  XORCY un1_inf_abs0_s_15 (
	.LI(un1_inf_abs0_axb_15),
	.CI(un1_inf_abs0_cry_14),
	.O(un1_inf_abs0_10[15])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_15_cZ (
	.DI(inf_abs0_2[15]),
	.CI(un1_inf_abs0_cry_14),
	.S(un1_inf_abs0_axb_15),
	.LO(un1_inf_abs0_cry_15)
);
// @7:74
  XORCY un1_inf_abs0_s_14 (
	.LI(un1_inf_abs0_axb_14),
	.CI(un1_inf_abs0_cry_13),
	.O(un1_inf_abs0_10[14])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_14_cZ (
	.DI(inf_abs0_2[14]),
	.CI(un1_inf_abs0_cry_13),
	.S(un1_inf_abs0_axb_14),
	.LO(un1_inf_abs0_cry_14)
);
// @7:74
  XORCY un1_inf_abs0_s_13 (
	.LI(un1_inf_abs0_axb_13),
	.CI(un1_inf_abs0_cry_12),
	.O(un1_inf_abs0_10[13])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_13_cZ (
	.DI(inf_abs0_2[13]),
	.CI(un1_inf_abs0_cry_12),
	.S(un1_inf_abs0_axb_13),
	.LO(un1_inf_abs0_cry_13)
);
// @7:74
  XORCY un1_inf_abs0_s_12 (
	.LI(un1_inf_abs0_axb_12),
	.CI(un1_inf_abs0_cry_11),
	.O(un1_inf_abs0_10[12])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_12_cZ (
	.DI(inf_abs0_2[12]),
	.CI(un1_inf_abs0_cry_11),
	.S(un1_inf_abs0_axb_12),
	.LO(un1_inf_abs0_cry_12)
);
// @7:74
  XORCY un1_inf_abs0_s_11 (
	.LI(un1_inf_abs0_axb_11),
	.CI(un1_inf_abs0_cry_10),
	.O(un1_inf_abs0_10[11])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_11_cZ (
	.DI(inf_abs0_2[11]),
	.CI(un1_inf_abs0_cry_10),
	.S(un1_inf_abs0_axb_11),
	.LO(un1_inf_abs0_cry_11)
);
// @7:74
  XORCY un1_inf_abs0_s_10 (
	.LI(un1_inf_abs0_axb_10),
	.CI(un1_inf_abs0_cry_9),
	.O(un1_inf_abs0_10[10])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_10_cZ (
	.DI(inf_abs0_2[10]),
	.CI(un1_inf_abs0_cry_9),
	.S(un1_inf_abs0_axb_10),
	.LO(un1_inf_abs0_cry_10)
);
// @7:74
  XORCY un1_inf_abs0_s_9 (
	.LI(un1_inf_abs0_axb_9),
	.CI(un1_inf_abs0_cry_8),
	.O(un1_inf_abs0_10[9])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_9_cZ (
	.DI(inf_abs0_2[9]),
	.CI(un1_inf_abs0_cry_8),
	.S(un1_inf_abs0_axb_9),
	.LO(un1_inf_abs0_cry_9)
);
// @7:74
  XORCY un1_inf_abs0_s_8 (
	.LI(un1_inf_abs0_axb_8),
	.CI(un1_inf_abs0_cry_7),
	.O(un1_inf_abs0_10[8])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_8_cZ (
	.DI(inf_abs0_2[8]),
	.CI(un1_inf_abs0_cry_7),
	.S(un1_inf_abs0_axb_8),
	.LO(un1_inf_abs0_cry_8)
);
// @7:74
  XORCY un1_inf_abs0_s_7 (
	.LI(un1_inf_abs0_axb_7),
	.CI(un1_inf_abs0_cry_6),
	.O(un1_inf_abs0_10[7])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_7_cZ (
	.DI(inf_abs0_2[7]),
	.CI(un1_inf_abs0_cry_6),
	.S(un1_inf_abs0_axb_7),
	.LO(un1_inf_abs0_cry_7)
);
// @7:74
  XORCY un1_inf_abs0_s_6 (
	.LI(un1_inf_abs0_axb_6),
	.CI(un1_inf_abs0_cry_5),
	.O(un1_inf_abs0_10[6])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_6_cZ (
	.DI(inf_abs0_2[6]),
	.CI(un1_inf_abs0_cry_5),
	.S(un1_inf_abs0_axb_6),
	.LO(un1_inf_abs0_cry_6)
);
// @7:74
  XORCY un1_inf_abs0_s_5 (
	.LI(un1_inf_abs0_axb_5),
	.CI(un1_inf_abs0_cry_4),
	.O(un1_inf_abs0_10[5])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_5_cZ (
	.DI(inf_abs0_2[5]),
	.CI(un1_inf_abs0_cry_4),
	.S(un1_inf_abs0_axb_5),
	.LO(un1_inf_abs0_cry_5)
);
// @7:74
  XORCY un1_inf_abs0_s_4 (
	.LI(un1_inf_abs0_axb_4),
	.CI(un1_inf_abs0_cry_3),
	.O(un1_inf_abs0_10[4])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_4_cZ (
	.DI(inf_abs0_2[4]),
	.CI(un1_inf_abs0_cry_3),
	.S(un1_inf_abs0_axb_4),
	.LO(un1_inf_abs0_cry_4)
);
// @7:74
  XORCY un1_inf_abs0_s_3 (
	.LI(un1_inf_abs0_axb_3),
	.CI(un1_inf_abs0_cry_2),
	.O(un1_inf_abs0_10[3])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_3_cZ (
	.DI(inf_abs0_2[3]),
	.CI(un1_inf_abs0_cry_2),
	.S(un1_inf_abs0_axb_3),
	.LO(un1_inf_abs0_cry_3)
);
// @7:74
  XORCY un1_inf_abs0_s_2 (
	.LI(un1_inf_abs0_axb_2),
	.CI(un1_inf_abs0_cry_1),
	.O(un1_inf_abs0_10[2])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_2_cZ (
	.DI(inf_abs0_2[2]),
	.CI(un1_inf_abs0_cry_1),
	.S(un1_inf_abs0_axb_2),
	.LO(un1_inf_abs0_cry_2)
);
// @7:74
  XORCY un1_inf_abs0_s_1 (
	.LI(un1_inf_abs0_axb_1),
	.CI(un1_inf_abs0_cry_0),
	.O(un1_inf_abs0_10[1])
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_1_cZ (
	.DI(inf_abs0_2[1]),
	.CI(un1_inf_abs0_cry_0),
	.S(un1_inf_abs0_axb_1),
	.LO(un1_inf_abs0_cry_1)
);
// @7:74
  MUXCY_L un1_inf_abs0_cry_0_cZ (
	.DI(inf_abs0_2[0]),
	.CI(GND),
	.S(un1_inf_abs0_10[0]),
	.LO(un1_inf_abs0_cry_0)
);
// @7:358
  XORCY un32_reg0_s_29_cZ (
	.LI(un32_reg0_axb_29),
	.CI(un32_reg0_cry_28),
	.O(un32_reg0_s_29)
);
// @7:358
  XORCY un32_reg0_s_28_cZ (
	.LI(un32_reg0_axb_28),
	.CI(un32_reg0_cry_27),
	.O(un32_reg0_s_28)
);
// @7:358
  MUXCY_L un32_reg0_cry_28_cZ (
	.DI(r_4[28]),
	.CI(un32_reg0_cry_27),
	.S(un32_reg0_axb_28),
	.LO(un32_reg0_cry_28)
);
// @7:358
  XORCY un32_reg0_s_27_cZ (
	.LI(un32_reg0_axb_27),
	.CI(un32_reg0_cry_26),
	.O(un32_reg0_s_27)
);
// @7:358
  MUXCY_L un32_reg0_cry_27_cZ (
	.DI(r_4[27]),
	.CI(un32_reg0_cry_26),
	.S(un32_reg0_axb_27),
	.LO(un32_reg0_cry_27)
);
// @7:358
  XORCY un32_reg0_s_26_cZ (
	.LI(un32_reg0_axb_26),
	.CI(un32_reg0_cry_25),
	.O(un32_reg0_s_26)
);
// @7:358
  MUXCY_L un32_reg0_cry_26_cZ (
	.DI(r_4[26]),
	.CI(un32_reg0_cry_25),
	.S(un32_reg0_axb_26),
	.LO(un32_reg0_cry_26)
);
// @7:358
  XORCY un32_reg0_s_25_cZ (
	.LI(un32_reg0_axb_25),
	.CI(un32_reg0_cry_24),
	.O(un32_reg0_s_25)
);
// @7:358
  MUXCY_L un32_reg0_cry_25_cZ (
	.DI(r_4[25]),
	.CI(un32_reg0_cry_24),
	.S(un32_reg0_axb_25),
	.LO(un32_reg0_cry_25)
);
// @7:358
  XORCY un32_reg0_s_24_cZ (
	.LI(un32_reg0_axb_24),
	.CI(un32_reg0_cry_23),
	.O(un32_reg0_s_24)
);
// @7:358
  MUXCY_L un32_reg0_cry_24_cZ (
	.DI(r_4[24]),
	.CI(un32_reg0_cry_23),
	.S(un32_reg0_axb_24),
	.LO(un32_reg0_cry_24)
);
// @7:358
  XORCY un32_reg0_s_23_cZ (
	.LI(un32_reg0_axb_23),
	.CI(un32_reg0_cry_22),
	.O(un32_reg0_s_23)
);
// @7:358
  MUXCY_L un32_reg0_cry_23_cZ (
	.DI(r_4[23]),
	.CI(un32_reg0_cry_22),
	.S(un32_reg0_axb_23),
	.LO(un32_reg0_cry_23)
);
// @7:358
  XORCY un32_reg0_s_22_cZ (
	.LI(un32_reg0_axb_22),
	.CI(un32_reg0_cry_21),
	.O(un32_reg0_s_22)
);
// @7:358
  MUXCY_L un32_reg0_cry_22_cZ (
	.DI(r_4[22]),
	.CI(un32_reg0_cry_21),
	.S(un32_reg0_axb_22),
	.LO(un32_reg0_cry_22)
);
// @7:358
  XORCY un32_reg0_s_21_cZ (
	.LI(un32_reg0_axb_21),
	.CI(un32_reg0_cry_20),
	.O(un32_reg0_s_21)
);
// @7:358
  MUXCY_L un32_reg0_cry_21_cZ (
	.DI(r_4[21]),
	.CI(un32_reg0_cry_20),
	.S(un32_reg0_axb_21),
	.LO(un32_reg0_cry_21)
);
// @7:358
  XORCY un32_reg0_s_20_cZ (
	.LI(un32_reg0_axb_20),
	.CI(un32_reg0_cry_19),
	.O(un32_reg0_s_20)
);
// @7:358
  MUXCY_L un32_reg0_cry_20_cZ (
	.DI(r_4[20]),
	.CI(un32_reg0_cry_19),
	.S(un32_reg0_axb_20),
	.LO(un32_reg0_cry_20)
);
// @7:358
  XORCY un32_reg0_s_19_cZ (
	.LI(un32_reg0_axb_19),
	.CI(un32_reg0_cry_18),
	.O(un32_reg0_s_19)
);
// @7:358
  MUXCY_L un32_reg0_cry_19_cZ (
	.DI(r_4[19]),
	.CI(un32_reg0_cry_18),
	.S(un32_reg0_axb_19),
	.LO(un32_reg0_cry_19)
);
// @7:358
  XORCY un32_reg0_s_18_cZ (
	.LI(un32_reg0_axb_18),
	.CI(un32_reg0_cry_17),
	.O(un32_reg0_s_18)
);
// @7:358
  MUXCY_L un32_reg0_cry_18_cZ (
	.DI(r_4[18]),
	.CI(un32_reg0_cry_17),
	.S(un32_reg0_axb_18),
	.LO(un32_reg0_cry_18)
);
// @7:358
  XORCY un32_reg0_s_17_cZ (
	.LI(un32_reg0_axb_17),
	.CI(un32_reg0_cry_16),
	.O(un32_reg0_s_17)
);
// @7:358
  MUXCY_L un32_reg0_cry_17_cZ (
	.DI(r_4[17]),
	.CI(un32_reg0_cry_16),
	.S(un32_reg0_axb_17),
	.LO(un32_reg0_cry_17)
);
// @7:358
  XORCY un32_reg0_s_16_cZ (
	.LI(un32_reg0_axb_16),
	.CI(un32_reg0_cry_15),
	.O(un32_reg0_s_16)
);
// @7:358
  MUXCY_L un32_reg0_cry_16_cZ (
	.DI(r_4[16]),
	.CI(un32_reg0_cry_15),
	.S(un32_reg0_axb_16),
	.LO(un32_reg0_cry_16)
);
// @7:358
  XORCY un32_reg0_s_15_cZ (
	.LI(un32_reg0_axb_15),
	.CI(un32_reg0_cry_14),
	.O(un32_reg0_s_15)
);
// @7:358
  MUXCY_L un32_reg0_cry_15_cZ (
	.DI(r_4[15]),
	.CI(un32_reg0_cry_14),
	.S(un32_reg0_axb_15),
	.LO(un32_reg0_cry_15)
);
// @7:358
  XORCY un32_reg0_s_14_cZ (
	.LI(un32_reg0_axb_14),
	.CI(un32_reg0_cry_13),
	.O(un32_reg0_s_14)
);
// @7:358
  MUXCY_L un32_reg0_cry_14_cZ (
	.DI(r_4[14]),
	.CI(un32_reg0_cry_13),
	.S(un32_reg0_axb_14),
	.LO(un32_reg0_cry_14)
);
// @7:358
  XORCY un32_reg0_s_13_cZ (
	.LI(un32_reg0_axb_13),
	.CI(un32_reg0_cry_12),
	.O(un32_reg0_s_13)
);
// @7:358
  MUXCY_L un32_reg0_cry_13_cZ (
	.DI(r_4[13]),
	.CI(un32_reg0_cry_12),
	.S(un32_reg0_axb_13),
	.LO(un32_reg0_cry_13)
);
// @7:358
  XORCY un32_reg0_s_12_cZ (
	.LI(un32_reg0_axb_12),
	.CI(un32_reg0_cry_11),
	.O(un32_reg0_s_12)
);
// @7:358
  MUXCY_L un32_reg0_cry_12_cZ (
	.DI(r_4[12]),
	.CI(un32_reg0_cry_11),
	.S(un32_reg0_axb_12),
	.LO(un32_reg0_cry_12)
);
// @7:358
  XORCY un32_reg0_s_11_cZ (
	.LI(un32_reg0_axb_11),
	.CI(un32_reg0_cry_10),
	.O(un32_reg0_s_11)
);
// @7:358
  MUXCY_L un32_reg0_cry_11_cZ (
	.DI(r_4[11]),
	.CI(un32_reg0_cry_10),
	.S(un32_reg0_axb_11),
	.LO(un32_reg0_cry_11)
);
// @7:358
  XORCY un32_reg0_s_10_cZ (
	.LI(un32_reg0_axb_10),
	.CI(un32_reg0_cry_9),
	.O(un32_reg0_s_10)
);
// @7:358
  MUXCY_L un32_reg0_cry_10_cZ (
	.DI(r_4[10]),
	.CI(un32_reg0_cry_9),
	.S(un32_reg0_axb_10),
	.LO(un32_reg0_cry_10)
);
// @7:358
  XORCY un32_reg0_s_9_cZ (
	.LI(un32_reg0_axb_9),
	.CI(un32_reg0_cry_8),
	.O(un32_reg0_s_9)
);
// @7:358
  MUXCY_L un32_reg0_cry_9_cZ (
	.DI(r_4[9]),
	.CI(un32_reg0_cry_8),
	.S(un32_reg0_axb_9),
	.LO(un32_reg0_cry_9)
);
// @7:358
  XORCY un32_reg0_s_8_cZ (
	.LI(un32_reg0_axb_8),
	.CI(un32_reg0_cry_7),
	.O(un32_reg0_s_8)
);
// @7:358
  MUXCY_L un32_reg0_cry_8_cZ (
	.DI(r_4[8]),
	.CI(un32_reg0_cry_7),
	.S(un32_reg0_axb_8),
	.LO(un32_reg0_cry_8)
);
// @7:358
  XORCY un32_reg0_s_7_cZ (
	.LI(un32_reg0_axb_7),
	.CI(un32_reg0_cry_6),
	.O(un32_reg0_s_7)
);
// @7:358
  MUXCY_L un32_reg0_cry_7_cZ (
	.DI(r_4[7]),
	.CI(un32_reg0_cry_6),
	.S(un32_reg0_axb_7),
	.LO(un32_reg0_cry_7)
);
// @7:358
  XORCY un32_reg0_s_6_cZ (
	.LI(un32_reg0_axb_6),
	.CI(un32_reg0_cry_5),
	.O(un32_reg0_s_6)
);
// @7:358
  MUXCY_L un32_reg0_cry_6_cZ (
	.DI(r_4[6]),
	.CI(un32_reg0_cry_5),
	.S(un32_reg0_axb_6),
	.LO(un32_reg0_cry_6)
);
// @7:358
  XORCY un32_reg0_s_5_cZ (
	.LI(un32_reg0_axb_5),
	.CI(un32_reg0_cry_4),
	.O(un32_reg0_s_5)
);
// @7:358
  MUXCY_L un32_reg0_cry_5_cZ (
	.DI(r_4[5]),
	.CI(un32_reg0_cry_4),
	.S(un32_reg0_axb_5),
	.LO(un32_reg0_cry_5)
);
// @7:358
  XORCY un32_reg0_s_4_cZ (
	.LI(un32_reg0_axb_4),
	.CI(un32_reg0_cry_3),
	.O(un32_reg0_s_4)
);
// @7:358
  MUXCY_L un32_reg0_cry_4_cZ (
	.DI(r_4[4]),
	.CI(un32_reg0_cry_3),
	.S(un32_reg0_axb_4),
	.LO(un32_reg0_cry_4)
);
// @7:358
  XORCY un32_reg0_s_3_cZ (
	.LI(un32_reg0_axb_3),
	.CI(un32_reg0_cry_2),
	.O(un32_reg0_s_3)
);
// @7:358
  MUXCY_L un32_reg0_cry_3_cZ (
	.DI(r_4[3]),
	.CI(un32_reg0_cry_2),
	.S(un32_reg0_axb_3),
	.LO(un32_reg0_cry_3)
);
// @7:358
  XORCY un32_reg0_s_2_cZ (
	.LI(un32_reg0_axb_2),
	.CI(un32_reg0_cry_1),
	.O(un32_reg0_s_2)
);
// @7:358
  MUXCY_L un32_reg0_cry_2_cZ (
	.DI(N_28),
	.CI(un32_reg0_cry_1),
	.S(un32_reg0_axb_2),
	.LO(un32_reg0_cry_2)
);
// @7:358
  XORCY un32_reg0_s_1_cZ (
	.LI(un32_reg0_axb_1),
	.CI(un32_reg0_cry_0),
	.O(un32_reg0_s_1)
);
// @7:358
  MUXCY_L un32_reg0_cry_1_cZ (
	.DI(r_4[1]),
	.CI(un32_reg0_cry_0),
	.S(un32_reg0_axb_1),
	.LO(un32_reg0_cry_1)
);
// @7:358
  MUXCY_L un32_reg0_cry_0_cZ (
	.DI(r_4[0]),
	.CI(VCC),
	.S(N_1035),
	.LO(un32_reg0_cry_0)
);
// @7:318
  XORCY un11_reg0_s_29_cZ (
	.LI(un11_reg0_axb_29),
	.CI(un11_reg0_cry_28),
	.O(un11_reg0_s_29)
);
// @7:318
  XORCY un11_reg0_s_28_cZ (
	.LI(un11_reg0_axb_28),
	.CI(un11_reg0_cry_27),
	.O(un11_reg0_s_28)
);
// @7:318
  MUXCY_L un11_reg0_cry_28_cZ (
	.DI(m_2[28]),
	.CI(un11_reg0_cry_27),
	.S(un11_reg0_axb_28),
	.LO(un11_reg0_cry_28)
);
// @7:318
  XORCY un11_reg0_s_27_cZ (
	.LI(un11_reg0_axb_27),
	.CI(un11_reg0_cry_26),
	.O(un11_reg0_s_27)
);
// @7:318
  MUXCY_L un11_reg0_cry_27_cZ (
	.DI(m_2[27]),
	.CI(un11_reg0_cry_26),
	.S(un11_reg0_axb_27),
	.LO(un11_reg0_cry_27)
);
// @7:318
  XORCY un11_reg0_s_26_cZ (
	.LI(un11_reg0_axb_26),
	.CI(un11_reg0_cry_25),
	.O(un11_reg0_s_26)
);
// @7:318
  MUXCY_L un11_reg0_cry_26_cZ (
	.DI(m_2[26]),
	.CI(un11_reg0_cry_25),
	.S(un11_reg0_axb_26),
	.LO(un11_reg0_cry_26)
);
// @7:318
  XORCY un11_reg0_s_25_cZ (
	.LI(un11_reg0_axb_25),
	.CI(un11_reg0_cry_24),
	.O(un11_reg0_s_25)
);
// @7:318
  MUXCY_L un11_reg0_cry_25_cZ (
	.DI(m_2[25]),
	.CI(un11_reg0_cry_24),
	.S(un11_reg0_axb_25),
	.LO(un11_reg0_cry_25)
);
// @7:318
  XORCY un11_reg0_s_24_cZ (
	.LI(un11_reg0_axb_24),
	.CI(un11_reg0_cry_23),
	.O(un11_reg0_s_24)
);
// @7:318
  MUXCY_L un11_reg0_cry_24_cZ (
	.DI(m_2[24]),
	.CI(un11_reg0_cry_23),
	.S(un11_reg0_axb_24),
	.LO(un11_reg0_cry_24)
);
// @7:318
  XORCY un11_reg0_s_23_cZ (
	.LI(un11_reg0_axb_23),
	.CI(un11_reg0_cry_22),
	.O(un11_reg0_s_23)
);
// @7:318
  MUXCY_L un11_reg0_cry_23_cZ (
	.DI(m_2[23]),
	.CI(un11_reg0_cry_22),
	.S(un11_reg0_axb_23),
	.LO(un11_reg0_cry_23)
);
// @7:318
  XORCY un11_reg0_s_22_cZ (
	.LI(un11_reg0_axb_22),
	.CI(un11_reg0_cry_21),
	.O(un11_reg0_s_22)
);
// @7:318
  MUXCY_L un11_reg0_cry_22_cZ (
	.DI(m_2[22]),
	.CI(un11_reg0_cry_21),
	.S(un11_reg0_axb_22),
	.LO(un11_reg0_cry_22)
);
// @7:318
  XORCY un11_reg0_s_21_cZ (
	.LI(un11_reg0_axb_21),
	.CI(un11_reg0_cry_20),
	.O(un11_reg0_s_21)
);
// @7:318
  MUXCY_L un11_reg0_cry_21_cZ (
	.DI(m_2[21]),
	.CI(un11_reg0_cry_20),
	.S(un11_reg0_axb_21),
	.LO(un11_reg0_cry_21)
);
// @7:318
  XORCY un11_reg0_s_20_cZ (
	.LI(un11_reg0_axb_20),
	.CI(un11_reg0_cry_19),
	.O(un11_reg0_s_20)
);
// @7:318
  MUXCY_L un11_reg0_cry_20_cZ (
	.DI(m_2[20]),
	.CI(un11_reg0_cry_19),
	.S(un11_reg0_axb_20),
	.LO(un11_reg0_cry_20)
);
// @7:318
  XORCY un11_reg0_s_19_cZ (
	.LI(un11_reg0_axb_19),
	.CI(un11_reg0_cry_18),
	.O(un11_reg0_s_19)
);
// @7:318
  MUXCY_L un11_reg0_cry_19_cZ (
	.DI(r_4[19]),
	.CI(un11_reg0_cry_18),
	.S(un11_reg0_axb_19),
	.LO(un11_reg0_cry_19)
);
// @7:318
  XORCY un11_reg0_s_18_cZ (
	.LI(un11_reg0_axb_18),
	.CI(un11_reg0_cry_17),
	.O(un11_reg0_s_18)
);
// @7:318
  MUXCY_L un11_reg0_cry_18_cZ (
	.DI(r_4[18]),
	.CI(un11_reg0_cry_17),
	.S(un11_reg0_axb_18),
	.LO(un11_reg0_cry_18)
);
// @7:318
  XORCY un11_reg0_s_17_cZ (
	.LI(un11_reg0_axb_17),
	.CI(un11_reg0_cry_16),
	.O(un11_reg0_s_17)
);
// @7:318
  MUXCY_L un11_reg0_cry_17_cZ (
	.DI(r_4[17]),
	.CI(un11_reg0_cry_16),
	.S(un11_reg0_axb_17),
	.LO(un11_reg0_cry_17)
);
// @7:318
  XORCY un11_reg0_s_16_cZ (
	.LI(un11_reg0_axb_16),
	.CI(un11_reg0_cry_15),
	.O(un11_reg0_s_16)
);
// @7:318
  MUXCY_L un11_reg0_cry_16_cZ (
	.DI(r_4[16]),
	.CI(un11_reg0_cry_15),
	.S(un11_reg0_axb_16),
	.LO(un11_reg0_cry_16)
);
// @7:318
  XORCY un11_reg0_s_15_cZ (
	.LI(un11_reg0_axb_15),
	.CI(un11_reg0_cry_14),
	.O(un11_reg0_s_15)
);
// @7:318
  MUXCY_L un11_reg0_cry_15_cZ (
	.DI(r_4[15]),
	.CI(un11_reg0_cry_14),
	.S(un11_reg0_axb_15),
	.LO(un11_reg0_cry_15)
);
// @7:318
  XORCY un11_reg0_s_14_cZ (
	.LI(un11_reg0_axb_14),
	.CI(un11_reg0_cry_13),
	.O(un11_reg0_s_14)
);
// @7:318
  MUXCY_L un11_reg0_cry_14_cZ (
	.DI(r_4[14]),
	.CI(un11_reg0_cry_13),
	.S(un11_reg0_axb_14),
	.LO(un11_reg0_cry_14)
);
// @7:318
  XORCY un11_reg0_s_13_cZ (
	.LI(un11_reg0_axb_13),
	.CI(un11_reg0_cry_12),
	.O(un11_reg0_s_13)
);
// @7:318
  MUXCY_L un11_reg0_cry_13_cZ (
	.DI(r_4[13]),
	.CI(un11_reg0_cry_12),
	.S(un11_reg0_axb_13),
	.LO(un11_reg0_cry_13)
);
// @7:318
  XORCY un11_reg0_s_12_cZ (
	.LI(un11_reg0_axb_12),
	.CI(un11_reg0_cry_11),
	.O(un11_reg0_s_12)
);
// @7:318
  MUXCY_L un11_reg0_cry_12_cZ (
	.DI(r_4[12]),
	.CI(un11_reg0_cry_11),
	.S(un11_reg0_axb_12),
	.LO(un11_reg0_cry_12)
);
// @7:318
  XORCY un11_reg0_s_11_cZ (
	.LI(un11_reg0_axb_11),
	.CI(un11_reg0_cry_10),
	.O(un11_reg0_s_11)
);
// @7:318
  MUXCY_L un11_reg0_cry_11_cZ (
	.DI(r_4[11]),
	.CI(un11_reg0_cry_10),
	.S(un11_reg0_axb_11),
	.LO(un11_reg0_cry_11)
);
// @7:318
  XORCY un11_reg0_s_10_cZ (
	.LI(un11_reg0_axb_10),
	.CI(un11_reg0_cry_9),
	.O(un11_reg0_s_10)
);
// @7:318
  MUXCY_L un11_reg0_cry_10_cZ (
	.DI(r_4[10]),
	.CI(un11_reg0_cry_9),
	.S(un11_reg0_axb_10),
	.LO(un11_reg0_cry_10)
);
// @7:318
  XORCY un11_reg0_s_9_cZ (
	.LI(un11_reg0_axb_9),
	.CI(un11_reg0_cry_8),
	.O(un11_reg0_s_9)
);
// @7:318
  MUXCY_L un11_reg0_cry_9_cZ (
	.DI(r_4[9]),
	.CI(un11_reg0_cry_8),
	.S(un11_reg0_axb_9),
	.LO(un11_reg0_cry_9)
);
// @7:318
  XORCY un11_reg0_s_8_cZ (
	.LI(un11_reg0_axb_8),
	.CI(un11_reg0_cry_7),
	.O(un11_reg0_s_8)
);
// @7:318
  MUXCY_L un11_reg0_cry_8_cZ (
	.DI(r_4[8]),
	.CI(un11_reg0_cry_7),
	.S(un11_reg0_axb_8),
	.LO(un11_reg0_cry_8)
);
// @7:318
  XORCY un11_reg0_s_7_cZ (
	.LI(un11_reg0_axb_7),
	.CI(un11_reg0_cry_6),
	.O(un11_reg0_s_7)
);
// @7:318
  MUXCY_L un11_reg0_cry_7_cZ (
	.DI(r_4[7]),
	.CI(un11_reg0_cry_6),
	.S(un11_reg0_axb_7),
	.LO(un11_reg0_cry_7)
);
// @7:318
  XORCY un11_reg0_s_6_cZ (
	.LI(un11_reg0_axb_6),
	.CI(un11_reg0_cry_5),
	.O(un11_reg0_s_6)
);
// @7:318
  MUXCY_L un11_reg0_cry_6_cZ (
	.DI(r_4[6]),
	.CI(un11_reg0_cry_5),
	.S(un11_reg0_axb_6),
	.LO(un11_reg0_cry_6)
);
// @7:318
  XORCY un11_reg0_s_5_cZ (
	.LI(un11_reg0_axb_5),
	.CI(un11_reg0_cry_4),
	.O(un11_reg0_s_5)
);
// @7:318
  MUXCY_L un11_reg0_cry_5_cZ (
	.DI(r_4[5]),
	.CI(un11_reg0_cry_4),
	.S(un11_reg0_axb_5),
	.LO(un11_reg0_cry_5)
);
// @7:318
  XORCY un11_reg0_s_4_cZ (
	.LI(un11_reg0_axb_4),
	.CI(un11_reg0_cry_3),
	.O(un11_reg0_s_4)
);
// @7:318
  MUXCY_L un11_reg0_cry_4_cZ (
	.DI(r_4[4]),
	.CI(un11_reg0_cry_3),
	.S(un11_reg0_axb_4),
	.LO(un11_reg0_cry_4)
);
// @7:318
  XORCY un11_reg0_s_3_cZ (
	.LI(un11_reg0_axb_3),
	.CI(un11_reg0_cry_2),
	.O(un11_reg0_s_3)
);
// @7:318
  MUXCY_L un11_reg0_cry_3_cZ (
	.DI(r_4[3]),
	.CI(un11_reg0_cry_2),
	.S(un11_reg0_axb_3),
	.LO(un11_reg0_cry_3)
);
// @7:318
  XORCY un11_reg0_s_2_cZ (
	.LI(un11_reg0_axb_2),
	.CI(un11_reg0_cry_1),
	.O(un11_reg0_s_2)
);
// @7:318
  MUXCY_L un11_reg0_cry_2_cZ (
	.DI(N_28),
	.CI(un11_reg0_cry_1),
	.S(un11_reg0_axb_2),
	.LO(un11_reg0_cry_2)
);
// @7:318
  XORCY un11_reg0_s_1_cZ (
	.LI(un11_reg0_axb_1),
	.CI(un11_reg0_cry_0),
	.O(un11_reg0_s_1)
);
// @7:318
  MUXCY_L un11_reg0_cry_1_cZ (
	.DI(r_4[1]),
	.CI(un11_reg0_cry_0),
	.S(un11_reg0_axb_1),
	.LO(un11_reg0_cry_1)
);
// @7:318
  MUXCY_L un11_reg0_cry_0_cZ (
	.DI(r_4[0]),
	.CI(GND),
	.S(un11_reg0_axb_0),
	.LO(un11_reg0_cry_0)
);
// @7:466
  XORCY un3_t_s_31_cZ (
	.LI(un3_t_axb_31),
	.CI(un3_t_cry_30),
	.O(un3_t_s_31)
);
// @7:466
  XORCY un3_t_s_30_cZ (
	.LI(un3_t_axb_30),
	.CI(un3_t_cry_29),
	.O(un3_t_s_30)
);
// @7:466
  MUXCY_L un3_t_cry_30_cZ (
	.DI(GND),
	.CI(un3_t_cry_29),
	.S(un3_t_axb_30),
	.LO(un3_t_cry_30)
);
// @7:466
  XORCY un3_t_s_29_cZ (
	.LI(un3_t_axb_29),
	.CI(un3_t_cry_28),
	.O(un3_t_s_29)
);
// @7:466
  MUXCY_L un3_t_cry_29_cZ (
	.DI(GND),
	.CI(un3_t_cry_28),
	.S(un3_t_axb_29),
	.LO(un3_t_cry_29)
);
// @7:466
  XORCY un3_t_s_28_cZ (
	.LI(un3_t_axb_28),
	.CI(un3_t_cry_27),
	.O(un3_t_s_28)
);
// @7:466
  MUXCY_L un3_t_cry_28_cZ (
	.DI(GND),
	.CI(un3_t_cry_27),
	.S(un3_t_axb_28),
	.LO(un3_t_cry_28)
);
// @7:466
  XORCY un3_t_s_27_cZ (
	.LI(un3_t_axb_27),
	.CI(un3_t_cry_26),
	.O(un3_t_s_27)
);
// @7:466
  MUXCY_L un3_t_cry_27_cZ (
	.DI(GND),
	.CI(un3_t_cry_26),
	.S(un3_t_axb_27),
	.LO(un3_t_cry_27)
);
// @7:466
  XORCY un3_t_s_26_cZ (
	.LI(un3_t_axb_26),
	.CI(un3_t_cry_25),
	.O(un3_t_s_26)
);
// @7:466
  MUXCY_L un3_t_cry_26_cZ (
	.DI(GND),
	.CI(un3_t_cry_25),
	.S(un3_t_axb_26),
	.LO(un3_t_cry_26)
);
// @7:466
  XORCY un3_t_s_25_cZ (
	.LI(un3_t_axb_25),
	.CI(un3_t_cry_24),
	.O(un3_t_s_25)
);
// @7:466
  MUXCY_L un3_t_cry_25_cZ (
	.DI(GND),
	.CI(un3_t_cry_24),
	.S(un3_t_axb_25),
	.LO(un3_t_cry_25)
);
// @7:466
  XORCY un3_t_s_24_cZ (
	.LI(un3_t_axb_24),
	.CI(un3_t_cry_23),
	.O(un3_t_s_24)
);
// @7:466
  MUXCY_L un3_t_cry_24_cZ (
	.DI(GND),
	.CI(un3_t_cry_23),
	.S(un3_t_axb_24),
	.LO(un3_t_cry_24)
);
// @7:466
  XORCY un3_t_s_23_cZ (
	.LI(un3_t_axb_23),
	.CI(un3_t_cry_22),
	.O(un3_t_s_23)
);
// @7:466
  MUXCY_L un3_t_cry_23_cZ (
	.DI(GND),
	.CI(un3_t_cry_22),
	.S(un3_t_axb_23),
	.LO(un3_t_cry_23)
);
// @7:466
  XORCY un3_t_s_22_cZ (
	.LI(un3_t_axb_22),
	.CI(un3_t_cry_21),
	.O(un3_t_s_22)
);
// @7:466
  MUXCY_L un3_t_cry_22_cZ (
	.DI(GND),
	.CI(un3_t_cry_21),
	.S(un3_t_axb_22),
	.LO(un3_t_cry_22)
);
// @7:466
  XORCY un3_t_s_21_cZ (
	.LI(un3_t_axb_21),
	.CI(un3_t_cry_20),
	.O(un3_t_s_21)
);
// @7:466
  MUXCY_L un3_t_cry_21_cZ (
	.DI(GND),
	.CI(un3_t_cry_20),
	.S(un3_t_axb_21),
	.LO(un3_t_cry_21)
);
// @7:466
  XORCY un3_t_s_20_cZ (
	.LI(un3_t_axb_20),
	.CI(un3_t_cry_19),
	.O(un3_t_s_20)
);
// @7:466
  MUXCY_L un3_t_cry_20_cZ (
	.DI(GND),
	.CI(un3_t_cry_19),
	.S(un3_t_axb_20),
	.LO(un3_t_cry_20)
);
// @7:466
  XORCY un3_t_s_19_cZ (
	.LI(un3_t_axb_19),
	.CI(un3_t_cry_18),
	.O(un3_t_s_19)
);
// @7:466
  MUXCY_L un3_t_cry_19_cZ (
	.DI(GND),
	.CI(un3_t_cry_18),
	.S(un3_t_axb_19),
	.LO(un3_t_cry_19)
);
// @7:466
  XORCY un3_t_s_18_cZ (
	.LI(un3_t_axb_18),
	.CI(un3_t_cry_17),
	.O(un3_t_s_18)
);
// @7:466
  MUXCY_L un3_t_cry_18_cZ (
	.DI(GND),
	.CI(un3_t_cry_17),
	.S(un3_t_axb_18),
	.LO(un3_t_cry_18)
);
// @7:466
  XORCY un3_t_s_17_cZ (
	.LI(un3_t_axb_17),
	.CI(un3_t_cry_16),
	.O(un3_t_s_17)
);
// @7:466
  MUXCY_L un3_t_cry_17_cZ (
	.DI(GND),
	.CI(un3_t_cry_16),
	.S(un3_t_axb_17),
	.LO(un3_t_cry_17)
);
// @7:466
  XORCY un3_t_s_16_cZ (
	.LI(un3_t_axb_16),
	.CI(un3_t_cry_15),
	.O(un3_t_s_16)
);
// @7:466
  MUXCY_L un3_t_cry_16_cZ (
	.DI(GND),
	.CI(un3_t_cry_15),
	.S(un3_t_axb_16),
	.LO(un3_t_cry_16)
);
// @7:466
  XORCY un3_t_s_15_cZ (
	.LI(un3_t_axb_15),
	.CI(un3_t_cry_14),
	.O(un3_t_s_15)
);
// @7:466
  MUXCY_L un3_t_cry_15_cZ (
	.DI(GND),
	.CI(un3_t_cry_14),
	.S(un3_t_axb_15),
	.LO(un3_t_cry_15)
);
// @7:466
  XORCY un3_t_s_14_cZ (
	.LI(un3_t_axb_14),
	.CI(un3_t_cry_13),
	.O(un3_t_s_14)
);
// @7:466
  MUXCY_L un3_t_cry_14_cZ (
	.DI(GND),
	.CI(un3_t_cry_13),
	.S(un3_t_axb_14),
	.LO(un3_t_cry_14)
);
// @7:466
  XORCY un3_t_s_13_cZ (
	.LI(un3_t_axb_13),
	.CI(un3_t_cry_12),
	.O(un3_t_s_13)
);
// @7:466
  MUXCY_L un3_t_cry_13_cZ (
	.DI(GND),
	.CI(un3_t_cry_12),
	.S(un3_t_axb_13),
	.LO(un3_t_cry_13)
);
// @7:466
  XORCY un3_t_s_12_cZ (
	.LI(un3_t_axb_12),
	.CI(un3_t_cry_11),
	.O(un3_t_s_12)
);
// @7:466
  MUXCY_L un3_t_cry_12_cZ (
	.DI(GND),
	.CI(un3_t_cry_11),
	.S(un3_t_axb_12),
	.LO(un3_t_cry_12)
);
// @7:466
  XORCY un3_t_s_11_cZ (
	.LI(un3_t_axb_11),
	.CI(un3_t_cry_10),
	.O(un3_t_s_11)
);
// @7:466
  MUXCY_L un3_t_cry_11_cZ (
	.DI(GND),
	.CI(un3_t_cry_10),
	.S(un3_t_axb_11),
	.LO(un3_t_cry_11)
);
// @7:466
  XORCY un3_t_s_10_cZ (
	.LI(un3_t_axb_10),
	.CI(un3_t_cry_9),
	.O(un3_t_s_10)
);
// @7:466
  MUXCY_L un3_t_cry_10_cZ (
	.DI(GND),
	.CI(un3_t_cry_9),
	.S(un3_t_axb_10),
	.LO(un3_t_cry_10)
);
// @7:466
  XORCY un3_t_s_9_cZ (
	.LI(un3_t_axb_9),
	.CI(un3_t_cry_8),
	.O(un3_t_s_9)
);
// @7:466
  MUXCY_L un3_t_cry_9_cZ (
	.DI(GND),
	.CI(un3_t_cry_8),
	.S(un3_t_axb_9),
	.LO(un3_t_cry_9)
);
// @7:466
  XORCY un3_t_s_8_cZ (
	.LI(un3_t_axb_8),
	.CI(un3_t_cry_7),
	.O(un3_t_s_8)
);
// @7:466
  MUXCY_L un3_t_cry_8_cZ (
	.DI(GND),
	.CI(un3_t_cry_7),
	.S(un3_t_axb_8),
	.LO(un3_t_cry_8)
);
// @7:466
  XORCY un3_t_s_7_cZ (
	.LI(un3_t_axb_7),
	.CI(un3_t_cry_6),
	.O(un3_t_s_7)
);
// @7:466
  MUXCY_L un3_t_cry_7_cZ (
	.DI(GND),
	.CI(un3_t_cry_6),
	.S(un3_t_axb_7),
	.LO(un3_t_cry_7)
);
// @7:466
  XORCY un3_t_s_6_cZ (
	.LI(un3_t_axb_6),
	.CI(un3_t_cry_5),
	.O(un3_t_s_6)
);
// @7:466
  MUXCY_L un3_t_cry_6_cZ (
	.DI(GND),
	.CI(un3_t_cry_5),
	.S(un3_t_axb_6),
	.LO(un3_t_cry_6)
);
// @7:466
  XORCY un3_t_s_5_cZ (
	.LI(un3_t_axb_5),
	.CI(un3_t_cry_4),
	.O(un3_t_s_5)
);
// @7:466
  MUXCY_L un3_t_cry_5_cZ (
	.DI(GND),
	.CI(un3_t_cry_4),
	.S(un3_t_axb_5),
	.LO(un3_t_cry_5)
);
// @7:466
  XORCY un3_t_s_4_cZ (
	.LI(un3_t_axb_4),
	.CI(un3_t_cry_3),
	.O(un3_t_s_4)
);
// @7:466
  MUXCY_L un3_t_cry_4_cZ (
	.DI(GND),
	.CI(un3_t_cry_3),
	.S(un3_t_axb_4),
	.LO(un3_t_cry_4)
);
// @7:466
  XORCY un3_t_s_3_cZ (
	.LI(un3_t_axb_3),
	.CI(un3_t_cry_2),
	.O(un3_t_s_3)
);
// @7:466
  MUXCY_L un3_t_cry_3_cZ (
	.DI(GND),
	.CI(un3_t_cry_2),
	.S(un3_t_axb_3),
	.LO(un3_t_cry_3)
);
// @7:466
  XORCY un3_t_s_2_cZ (
	.LI(un3_t_axb_2),
	.CI(un3_t_cry_1),
	.O(un3_t_s_2)
);
// @7:466
  MUXCY_L un3_t_cry_2_cZ (
	.DI(GND),
	.CI(un3_t_cry_1),
	.S(un3_t_axb_2),
	.LO(un3_t_cry_2)
);
// @7:466
  XORCY un3_t_s_1_cZ (
	.LI(un3_t_axb_1),
	.CI(un3_t_cry_0),
	.O(un3_t_s_1)
);
// @7:466
  MUXCY_L un3_t_cry_1_cZ (
	.DI(GND),
	.CI(un3_t_cry_0),
	.S(un3_t_axb_1),
	.LO(un3_t_cry_1)
);
// @7:466
  MUXCY_L un3_t_cry_0_cZ (
	.DI(GND),
	.CI(un3_t_cry_0_cy),
	.S(un3_t_axb_0),
	.LO(un3_t_cry_0)
);
// @7:243
  XORCY reg3_1_1_s_31 (
	.LI(reg3_1_1_axb_31),
	.CI(reg3_1_1_cry_30),
	.O(reg3_1_1[31])
);
// @7:243
  XORCY reg3_1_1_s_30 (
	.LI(reg3_1_1_axb_30),
	.CI(reg3_1_1_cry_29),
	.O(reg3_1_1[30])
);
// @7:243
  MUXCY_L reg3_1_1_cry_30_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_29),
	.S(reg3_1_1_axb_30),
	.LO(reg3_1_1_cry_30)
);
// @7:243
  XORCY reg3_1_1_s_29 (
	.LI(reg3_1_1_axb_29),
	.CI(reg3_1_1_cry_28),
	.O(reg3_1_1[29])
);
// @7:243
  MUXCY_L reg3_1_1_cry_29_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_28),
	.S(reg3_1_1_axb_29),
	.LO(reg3_1_1_cry_29)
);
// @7:243
  XORCY reg3_1_1_s_28 (
	.LI(reg3_1_1_axb_28),
	.CI(reg3_1_1_cry_27),
	.O(reg3_1_1[28])
);
// @7:243
  MUXCY_L reg3_1_1_cry_28_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_27),
	.S(reg3_1_1_axb_28),
	.LO(reg3_1_1_cry_28)
);
// @7:243
  XORCY reg3_1_1_s_27 (
	.LI(reg3_1_1_axb_27),
	.CI(reg3_1_1_cry_26),
	.O(reg3_1_1[27])
);
// @7:243
  MUXCY_L reg3_1_1_cry_27_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_26),
	.S(reg3_1_1_axb_27),
	.LO(reg3_1_1_cry_27)
);
// @7:243
  XORCY reg3_1_1_s_26 (
	.LI(reg3_1_1_axb_26),
	.CI(reg3_1_1_cry_25),
	.O(reg3_1_1[26])
);
// @7:243
  MUXCY_L reg3_1_1_cry_26_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_25),
	.S(reg3_1_1_axb_26),
	.LO(reg3_1_1_cry_26)
);
// @7:243
  XORCY reg3_1_1_s_25 (
	.LI(reg3_1_1_axb_25),
	.CI(reg3_1_1_cry_24),
	.O(reg3_1_1[25])
);
// @7:243
  MUXCY_L reg3_1_1_cry_25_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_24),
	.S(reg3_1_1_axb_25),
	.LO(reg3_1_1_cry_25)
);
// @7:243
  XORCY reg3_1_1_s_24 (
	.LI(reg3_1_1_axb_24),
	.CI(reg3_1_1_cry_23),
	.O(reg3_1_1[24])
);
// @7:243
  MUXCY_L reg3_1_1_cry_24_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_23),
	.S(reg3_1_1_axb_24),
	.LO(reg3_1_1_cry_24)
);
// @7:243
  XORCY reg3_1_1_s_23 (
	.LI(reg3_1_1_axb_23),
	.CI(reg3_1_1_cry_22),
	.O(reg3_1_1[23])
);
// @7:243
  MUXCY_L reg3_1_1_cry_23_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_22),
	.S(reg3_1_1_axb_23),
	.LO(reg3_1_1_cry_23)
);
// @7:243
  XORCY reg3_1_1_s_22 (
	.LI(reg3_1_1_axb_22),
	.CI(reg3_1_1_cry_21),
	.O(reg3_1_1[22])
);
// @7:243
  MUXCY_L reg3_1_1_cry_22_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_21),
	.S(reg3_1_1_axb_22),
	.LO(reg3_1_1_cry_22)
);
// @7:243
  XORCY reg3_1_1_s_21 (
	.LI(reg3_1_1_axb_21),
	.CI(reg3_1_1_cry_20),
	.O(reg3_1_1[21])
);
// @7:243
  MUXCY_L reg3_1_1_cry_21_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_20),
	.S(reg3_1_1_axb_21),
	.LO(reg3_1_1_cry_21)
);
// @7:243
  XORCY reg3_1_1_s_20 (
	.LI(reg3_1_1_axb_20),
	.CI(reg3_1_1_cry_19),
	.O(reg3_1_1[20])
);
// @7:243
  MUXCY_L reg3_1_1_cry_20_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_19),
	.S(reg3_1_1_axb_20),
	.LO(reg3_1_1_cry_20)
);
// @7:243
  XORCY reg3_1_1_s_19 (
	.LI(reg3_1_1_axb_19),
	.CI(reg3_1_1_cry_18),
	.O(reg3_1_1[19])
);
// @7:243
  MUXCY_L reg3_1_1_cry_19_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_18),
	.S(reg3_1_1_axb_19),
	.LO(reg3_1_1_cry_19)
);
// @7:243
  XORCY reg3_1_1_s_18 (
	.LI(reg3_1_1_axb_18),
	.CI(reg3_1_1_cry_17),
	.O(reg3_1_1[18])
);
// @7:243
  MUXCY_L reg3_1_1_cry_18_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_17),
	.S(reg3_1_1_axb_18),
	.LO(reg3_1_1_cry_18)
);
// @7:243
  XORCY reg3_1_1_s_17 (
	.LI(reg3_1_1_axb_17),
	.CI(reg3_1_1_cry_16),
	.O(reg3_1_1[17])
);
// @7:243
  MUXCY_L reg3_1_1_cry_17_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_16),
	.S(reg3_1_1_axb_17),
	.LO(reg3_1_1_cry_17)
);
// @7:243
  XORCY reg3_1_1_s_16 (
	.LI(reg3_1_1_axb_16),
	.CI(reg3_1_1_cry_15),
	.O(reg3_1_1[16])
);
// @7:243
  MUXCY_L reg3_1_1_cry_16_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_15),
	.S(reg3_1_1_axb_16),
	.LO(reg3_1_1_cry_16)
);
// @7:243
  XORCY reg3_1_1_s_15 (
	.LI(reg3_1_1_axb_15),
	.CI(reg3_1_1_cry_14),
	.O(reg3_1_1[15])
);
// @7:243
  MUXCY_L reg3_1_1_cry_15_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_14),
	.S(reg3_1_1_axb_15),
	.LO(reg3_1_1_cry_15)
);
// @7:243
  XORCY reg3_1_1_s_14 (
	.LI(reg3_1_1_axb_14),
	.CI(reg3_1_1_cry_13),
	.O(reg3_1_1[14])
);
// @7:243
  MUXCY_L reg3_1_1_cry_14_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_13),
	.S(reg3_1_1_axb_14),
	.LO(reg3_1_1_cry_14)
);
// @7:243
  XORCY reg3_1_1_s_13 (
	.LI(reg3_1_1_axb_13),
	.CI(reg3_1_1_cry_12),
	.O(reg3_1_1[13])
);
// @7:243
  MUXCY_L reg3_1_1_cry_13_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_12),
	.S(reg3_1_1_axb_13),
	.LO(reg3_1_1_cry_13)
);
// @7:243
  XORCY reg3_1_1_s_12 (
	.LI(reg3_1_1_axb_12),
	.CI(reg3_1_1_cry_11),
	.O(reg3_1_1[12])
);
// @7:243
  MUXCY_L reg3_1_1_cry_12_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_11),
	.S(reg3_1_1_axb_12),
	.LO(reg3_1_1_cry_12)
);
// @7:243
  XORCY reg3_1_1_s_11 (
	.LI(reg3_1_1_axb_11),
	.CI(reg3_1_1_cry_10),
	.O(reg3_1_1[11])
);
// @7:243
  MUXCY_L reg3_1_1_cry_11_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_10),
	.S(reg3_1_1_axb_11),
	.LO(reg3_1_1_cry_11)
);
// @7:243
  XORCY reg3_1_1_s_10 (
	.LI(reg3_1_1_axb_10),
	.CI(reg3_1_1_cry_9),
	.O(reg3_1_1[10])
);
// @7:243
  MUXCY_L reg3_1_1_cry_10_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_9),
	.S(reg3_1_1_axb_10),
	.LO(reg3_1_1_cry_10)
);
// @7:243
  XORCY reg3_1_1_s_9 (
	.LI(reg3_1_1_axb_9),
	.CI(reg3_1_1_cry_8),
	.O(reg3_1_1[9])
);
// @7:243
  MUXCY_L reg3_1_1_cry_9_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_8),
	.S(reg3_1_1_axb_9),
	.LO(reg3_1_1_cry_9)
);
// @7:243
  XORCY reg3_1_1_s_8 (
	.LI(reg3_1_1_axb_8),
	.CI(reg3_1_1_cry_7),
	.O(reg3_1_1[8])
);
// @7:243
  MUXCY_L reg3_1_1_cry_8_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_7),
	.S(reg3_1_1_axb_8),
	.LO(reg3_1_1_cry_8)
);
// @7:243
  XORCY reg3_1_1_s_7 (
	.LI(reg3_1_1_axb_7),
	.CI(reg3_1_1_cry_6),
	.O(reg3_1_1[7])
);
// @7:243
  MUXCY_L reg3_1_1_cry_7_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_6),
	.S(reg3_1_1_axb_7),
	.LO(reg3_1_1_cry_7)
);
// @7:243
  XORCY reg3_1_1_s_6 (
	.LI(reg3_1_1_axb_6),
	.CI(reg3_1_1_cry_5),
	.O(reg3_1_1[6])
);
// @7:243
  MUXCY_L reg3_1_1_cry_6_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_5),
	.S(reg3_1_1_axb_6),
	.LO(reg3_1_1_cry_6)
);
// @7:243
  XORCY reg3_1_1_s_5 (
	.LI(reg3_1_1_axb_5),
	.CI(reg3_1_1_cry_4),
	.O(reg3_1_1[5])
);
// @7:243
  MUXCY_L reg3_1_1_cry_5_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_4),
	.S(reg3_1_1_axb_5),
	.LO(reg3_1_1_cry_5)
);
// @7:243
  XORCY reg3_1_1_s_4 (
	.LI(reg3_1_1_axb_4),
	.CI(reg3_1_1_cry_3),
	.O(reg3_1_1[4])
);
// @7:243
  MUXCY_L reg3_1_1_cry_4_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_3),
	.S(reg3_1_1_axb_4),
	.LO(reg3_1_1_cry_4)
);
// @7:243
  XORCY reg3_1_1_s_3 (
	.LI(reg3_1_1_axb_3),
	.CI(reg3_1_1_cry_2),
	.O(reg3_1_1[3])
);
// @7:243
  MUXCY_L reg3_1_1_cry_3_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_2),
	.S(reg3_1_1_axb_3),
	.LO(reg3_1_1_cry_3)
);
// @7:243
  XORCY reg3_1_1_s_2 (
	.LI(reg3_1_1_axb_2),
	.CI(reg3_1_1_cry_1),
	.O(reg3_1_1[2])
);
// @7:243
  MUXCY_L reg3_1_1_cry_2_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_1),
	.S(reg3_1_1_axb_2),
	.LO(reg3_1_1_cry_2)
);
// @7:243
  XORCY reg3_1_1_s_1 (
	.LI(reg3_1_1_axb_1),
	.CI(reg3_1_1_cry_0),
	.O(reg3_1_1[1])
);
// @7:243
  MUXCY_L reg3_1_1_cry_1_cZ (
	.DI(GND),
	.CI(reg3_1_1_cry_0),
	.S(reg3_1_1_axb_1),
	.LO(reg3_1_1_cry_1)
);
// @7:243
  MUXCY_L reg3_1_1_cry_0_cZ (
	.DI(GND),
	.CI(VCC),
	.S(reg3_1_1_axb_0),
	.LO(reg3_1_1_cry_0)
);
// @7:83
  XORCY inf_abs0_2_s_30 (
	.LI(inf_abs0_2_axb_30),
	.CI(inf_abs0_2_cry_29),
	.O(inf_abs0_2[30])
);
// @7:83
  MUXCY inf_abs0_2_cry_30 (
	.DI(GND),
	.CI(inf_abs0_2_cry_29),
	.S(inf_abs0_2_axb_30),
	.O(inf_abs0_2_0[31])
);
// @7:83
  XORCY inf_abs0_2_s_29 (
	.LI(inf_abs0_2_axb_29),
	.CI(inf_abs0_2_cry_28),
	.O(inf_abs0_2[29])
);
// @7:83
  XORCY inf_abs0_2_s_28 (
	.LI(inf_abs0_2_axb_28),
	.CI(inf_abs0_2_cry_27),
	.O(inf_abs0_2[28])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_28_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_27),
	.S(inf_abs0_2_axb_28),
	.LO(inf_abs0_2_cry_28)
);
// @7:83
  XORCY inf_abs0_2_s_27 (
	.LI(inf_abs0_2_axb_27),
	.CI(inf_abs0_2_cry_26),
	.O(inf_abs0_2[27])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_27_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_26),
	.S(inf_abs0_2_axb_27),
	.LO(inf_abs0_2_cry_27)
);
// @7:83
  XORCY inf_abs0_2_s_26 (
	.LI(inf_abs0_2_axb_26),
	.CI(inf_abs0_2_cry_25),
	.O(inf_abs0_2[26])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_26_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_25),
	.S(inf_abs0_2_axb_26),
	.LO(inf_abs0_2_cry_26)
);
// @7:83
  XORCY inf_abs0_2_s_25 (
	.LI(inf_abs0_2_axb_25),
	.CI(inf_abs0_2_cry_24),
	.O(inf_abs0_2[25])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_25_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_24),
	.S(inf_abs0_2_axb_25),
	.LO(inf_abs0_2_cry_25)
);
// @7:83
  XORCY inf_abs0_2_s_24 (
	.LI(inf_abs0_2_axb_24),
	.CI(inf_abs0_2_cry_23),
	.O(inf_abs0_2[24])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_24_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_23),
	.S(inf_abs0_2_axb_24),
	.LO(inf_abs0_2_cry_24)
);
// @7:83
  XORCY inf_abs0_2_s_23 (
	.LI(inf_abs0_2_axb_23),
	.CI(inf_abs0_2_cry_22),
	.O(inf_abs0_2[23])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_23_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_22),
	.S(inf_abs0_2_axb_23),
	.LO(inf_abs0_2_cry_23)
);
// @7:83
  XORCY inf_abs0_2_s_22 (
	.LI(inf_abs0_2_axb_22),
	.CI(inf_abs0_2_cry_21),
	.O(inf_abs0_2[22])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_22_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_21),
	.S(inf_abs0_2_axb_22),
	.LO(inf_abs0_2_cry_22)
);
// @7:83
  XORCY inf_abs0_2_s_21 (
	.LI(inf_abs0_2_axb_21),
	.CI(inf_abs0_2_cry_20),
	.O(inf_abs0_2[21])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_21_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_20),
	.S(inf_abs0_2_axb_21),
	.LO(inf_abs0_2_cry_21)
);
// @7:83
  XORCY inf_abs0_2_s_20 (
	.LI(inf_abs0_2_axb_20),
	.CI(inf_abs0_2_cry_19),
	.O(inf_abs0_2[20])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_20_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_19),
	.S(inf_abs0_2_axb_20),
	.LO(inf_abs0_2_cry_20)
);
// @7:83
  XORCY inf_abs0_2_s_19 (
	.LI(inf_abs0_2_axb_19),
	.CI(inf_abs0_2_cry_18),
	.O(inf_abs0_2[19])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_19_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_18),
	.S(inf_abs0_2_axb_19),
	.LO(inf_abs0_2_cry_19)
);
// @7:83
  XORCY inf_abs0_2_s_18 (
	.LI(inf_abs0_2_axb_18),
	.CI(inf_abs0_2_cry_17),
	.O(inf_abs0_2[18])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_18_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_17),
	.S(inf_abs0_2_axb_18),
	.LO(inf_abs0_2_cry_18)
);
// @7:83
  XORCY inf_abs0_2_s_17 (
	.LI(inf_abs0_2_axb_17),
	.CI(inf_abs0_2_cry_16),
	.O(inf_abs0_2[17])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_17_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_16),
	.S(inf_abs0_2_axb_17),
	.LO(inf_abs0_2_cry_17)
);
// @7:83
  XORCY inf_abs0_2_s_16 (
	.LI(inf_abs0_2_axb_16),
	.CI(inf_abs0_2_cry_15),
	.O(inf_abs0_2[16])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_16_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_15),
	.S(inf_abs0_2_axb_16),
	.LO(inf_abs0_2_cry_16)
);
// @7:83
  XORCY inf_abs0_2_s_15 (
	.LI(inf_abs0_2_axb_15),
	.CI(inf_abs0_2_cry_14),
	.O(inf_abs0_2[15])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_15_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_14),
	.S(inf_abs0_2_axb_15),
	.LO(inf_abs0_2_cry_15)
);
// @7:83
  XORCY inf_abs0_2_s_14 (
	.LI(inf_abs0_2_axb_14),
	.CI(inf_abs0_2_cry_13),
	.O(inf_abs0_2[14])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_14_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_13),
	.S(inf_abs0_2_axb_14),
	.LO(inf_abs0_2_cry_14)
);
// @7:83
  XORCY inf_abs0_2_s_13 (
	.LI(inf_abs0_2_axb_13),
	.CI(inf_abs0_2_cry_12),
	.O(inf_abs0_2[13])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_13_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_12),
	.S(inf_abs0_2_axb_13),
	.LO(inf_abs0_2_cry_13)
);
// @7:83
  XORCY inf_abs0_2_s_12 (
	.LI(inf_abs0_2_axb_12),
	.CI(inf_abs0_2_cry_11),
	.O(inf_abs0_2[12])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_12_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_11),
	.S(inf_abs0_2_axb_12),
	.LO(inf_abs0_2_cry_12)
);
// @7:83
  XORCY inf_abs0_2_s_11 (
	.LI(inf_abs0_2_axb_11),
	.CI(inf_abs0_2_cry_10),
	.O(inf_abs0_2[11])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_11_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_10),
	.S(inf_abs0_2_axb_11),
	.LO(inf_abs0_2_cry_11)
);
// @7:83
  XORCY inf_abs0_2_s_10 (
	.LI(inf_abs0_2_axb_10),
	.CI(inf_abs0_2_cry_9),
	.O(inf_abs0_2[10])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_10_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_9),
	.S(inf_abs0_2_axb_10),
	.LO(inf_abs0_2_cry_10)
);
// @7:83
  XORCY inf_abs0_2_s_9 (
	.LI(inf_abs0_2_axb_9),
	.CI(inf_abs0_2_cry_8),
	.O(inf_abs0_2[9])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_9_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_8),
	.S(inf_abs0_2_axb_9),
	.LO(inf_abs0_2_cry_9)
);
// @7:83
  XORCY inf_abs0_2_s_8 (
	.LI(inf_abs0_2_axb_8),
	.CI(inf_abs0_2_cry_7),
	.O(inf_abs0_2[8])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_8_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_7),
	.S(inf_abs0_2_axb_8),
	.LO(inf_abs0_2_cry_8)
);
// @7:83
  XORCY inf_abs0_2_s_7 (
	.LI(inf_abs0_2_axb_7),
	.CI(inf_abs0_2_cry_6),
	.O(inf_abs0_2[7])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_7_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_6),
	.S(inf_abs0_2_axb_7),
	.LO(inf_abs0_2_cry_7)
);
// @7:83
  XORCY inf_abs0_2_s_6 (
	.LI(inf_abs0_2_axb_6),
	.CI(inf_abs0_2_cry_5),
	.O(inf_abs0_2[6])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_6_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_5),
	.S(inf_abs0_2_axb_6),
	.LO(inf_abs0_2_cry_6)
);
// @7:83
  XORCY inf_abs0_2_s_5 (
	.LI(inf_abs0_2_axb_5),
	.CI(inf_abs0_2_cry_4),
	.O(inf_abs0_2[5])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_5_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_4),
	.S(inf_abs0_2_axb_5),
	.LO(inf_abs0_2_cry_5)
);
// @7:83
  XORCY inf_abs0_2_s_4 (
	.LI(inf_abs0_2_axb_4),
	.CI(inf_abs0_2_cry_3),
	.O(inf_abs0_2[4])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_4_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_3),
	.S(inf_abs0_2_axb_4),
	.LO(inf_abs0_2_cry_4)
);
// @7:83
  XORCY inf_abs0_2_s_3 (
	.LI(inf_abs0_2_axb_3),
	.CI(inf_abs0_2_cry_2),
	.O(inf_abs0_2[3])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_3_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_2),
	.S(inf_abs0_2_axb_3),
	.LO(inf_abs0_2_cry_3)
);
// @7:83
  XORCY inf_abs0_2_s_2 (
	.LI(inf_abs0_2_axb_2),
	.CI(inf_abs0_2_cry_1),
	.O(inf_abs0_2[2])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_2_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_1),
	.S(inf_abs0_2_axb_2),
	.LO(inf_abs0_2_cry_2)
);
// @7:83
  XORCY inf_abs0_2_s_1 (
	.LI(inf_abs0_2_axb_1),
	.CI(inf_abs0_2_cry_0),
	.O(inf_abs0_2[1])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_1_cZ (
	.DI(GND),
	.CI(inf_abs0_2_cry_0),
	.S(inf_abs0_2_axb_1),
	.LO(inf_abs0_2_cry_1)
);
// @7:83
  XORCY inf_abs0_2_s_0 (
	.LI(inf_abs0_2_axb_0),
	.CI(ir_fast[31]),
	.O(inf_abs0_2[0])
);
// @7:83
  MUXCY_L inf_abs0_2_cry_0_cZ (
	.DI(GND),
	.CI(ir_fast[31]),
	.S(inf_abs0_2_axb_0),
	.LO(inf_abs0_2_cry_0)
);
// @7:151
  LUT4 un26_r_lt30_cZ (
	.I0(m_2_i[31]),
	.I1(m_2[30]),
	.I2(r_4_i[31]),
	.I3(r_6[30]),
	.O(un26_r_lt30)
);
defparam un26_r_lt30_cZ.INIT=16'h0A8E;
// @7:151
  MUXCY_L \un26_r_cry_cZ[28]  (
	.DI(un26_r_lt28),
	.CI(un26_r_cry[26]),
	.S(un26_r_df28),
	.LO(un26_r_cry[28])
);
// @7:151
  MUXCY_L \un26_r_cry_cZ[26]  (
	.DI(un26_r_lt26),
	.CI(un26_r_cry[24]),
	.S(un26_r_df26),
	.LO(un26_r_cry[26])
);
// @7:151
  MUXCY_L \un26_r_cry_cZ[24]  (
	.DI(un26_r_lt24),
	.CI(un26_r_cry[22]),
	.S(un26_r_df24),
	.LO(un26_r_cry[24])
);
// @7:151
  MUXCY_L \un26_r_cry_cZ[22]  (
	.DI(un26_r_lt22),
	.CI(un26_r_cry[20]),
	.S(un26_r_df22),
	.LO(un26_r_cry[22])
);
// @7:151
  MUXCY_L \un26_r_cry_cZ[20]  (
	.DI(un26_r_lt20),
	.CI(un26_r_cry[18]),
	.S(un26_r_df20),
	.LO(un26_r_cry[20])
);
// @7:151
  MUXCY_L \un26_r_cry_cZ[18]  (
	.DI(un26_r_lt18),
	.CI(un26_r_cry[16]),
	.S(un26_r_df18),
	.LO(un26_r_cry[18])
);
// @7:151
  LUT4 un26_r_lt18_cZ (
	.I0(m_2[19]),
	.I1(m_2[18]),
	.I2(r_4[19]),
	.I3(r_4[18]),
	.O(un26_r_lt18)
);
defparam un26_r_lt18_cZ.INIT=16'h0A8E;
// @7:151
  MUXCY_L \un26_r_cry_cZ[16]  (
	.DI(un26_r_lt16),
	.CI(un26_r_cry[14]),
	.S(un26_r_df16),
	.LO(un26_r_cry[16])
);
// @7:151
  LUT4 un26_r_lt16_cZ (
	.I0(m_2[16]),
	.I1(m_2[17]),
	.I2(r_4[16]),
	.I3(r_4[17]),
	.O(un26_r_lt16)
);
defparam un26_r_lt16_cZ.INIT=16'h08CE;
// @7:151
  MUXCY_L \un26_r_cry_cZ[14]  (
	.DI(un26_r_lt14),
	.CI(un26_r_cry[12]),
	.S(un26_r_df14),
	.LO(un26_r_cry[14])
);
// @7:151
  LUT4 un26_r_lt14_cZ (
	.I0(m_2[14]),
	.I1(m_2[15]),
	.I2(r_4[14]),
	.I3(r_4[15]),
	.O(un26_r_lt14)
);
defparam un26_r_lt14_cZ.INIT=16'h08CE;
// @7:151
  MUXCY_L \un26_r_cry_cZ[12]  (
	.DI(un26_r_lt12),
	.CI(un26_r_cry[10]),
	.S(un26_r_df12),
	.LO(un26_r_cry[12])
);
// @7:151
  LUT4 un26_r_lt12_cZ (
	.I0(m_2[12]),
	.I1(m_2[13]),
	.I2(r_4[12]),
	.I3(r_4[13]),
	.O(un26_r_lt12)
);
defparam un26_r_lt12_cZ.INIT=16'h08CE;
// @7:151
  MUXCY_L \un26_r_cry_cZ[10]  (
	.DI(un26_r_lt10),
	.CI(un26_r_cry[8]),
	.S(un26_r_df10),
	.LO(un26_r_cry[10])
);
// @7:151
  LUT4 un26_r_lt10_cZ (
	.I0(m_2[10]),
	.I1(m_2[11]),
	.I2(r_4[11]),
	.I3(r_4[10]),
	.O(un26_r_lt10)
);
defparam un26_r_lt10_cZ.INIT=16'h0C8E;
// @7:151
  MUXCY_L \un26_r_cry_cZ[8]  (
	.DI(un26_r_lt8),
	.CI(un26_r_cry[6]),
	.S(un26_r_df8),
	.LO(un26_r_cry[8])
);
// @7:151
  LUT4 un26_r_lt8_cZ (
	.I0(m_2[8]),
	.I1(m_2[9]),
	.I2(r_4[8]),
	.I3(r_4[9]),
	.O(un26_r_lt8)
);
defparam un26_r_lt8_cZ.INIT=16'h08CE;
// @7:151
  MUXCY_L \un26_r_cry_cZ[6]  (
	.DI(un26_r_lt6),
	.CI(un26_r_cry[4]),
	.S(un26_r_df6),
	.LO(un26_r_cry[6])
);
// @7:151
  LUT4 un26_r_lt6_cZ (
	.I0(m_2[7]),
	.I1(m_2[6]),
	.I2(r_4[6]),
	.I3(r_4[7]),
	.O(un26_r_lt6)
);
defparam un26_r_lt6_cZ.INIT=16'h08AE;
// @7:151
  MUXCY_L \un26_r_cry_cZ[4]  (
	.DI(un26_r_lt4),
	.CI(un26_r_cry[2]),
	.S(un26_r_df4),
	.LO(un26_r_cry[4])
);
// @7:151
  LUT4 un26_r_lt4_cZ (
	.I0(m_2[4]),
	.I1(m_2[5]),
	.I2(r_4[4]),
	.I3(r_4[5]),
	.O(un26_r_lt4)
);
defparam un26_r_lt4_cZ.INIT=16'h08CE;
// @7:151
  MUXCY_L \un26_r_cry_cZ[2]  (
	.DI(un26_r_lt2),
	.CI(un26_r_cry[0]),
	.S(un26_r_df2),
	.LO(un26_r_cry[2])
);
// @7:151
  LUT4 un26_r_lt2_cZ (
	.I0(m_2[2]),
	.I1(m_2[3]),
	.I2(r_4[3]),
	.I3(N_28),
	.O(un26_r_lt2)
);
defparam un26_r_lt2_cZ.INIT=16'h0C8E;
// @7:151
  MUXCY_L \un26_r_cry_cZ[0]  (
	.DI(un26_r_lt0),
	.CI(GND),
	.S(un26_r_df0),
	.LO(un26_r_cry[0])
);
// @7:151
  LUT4 un26_r_lt0_cZ (
	.I0(m_2[1]),
	.I1(m_2[0]),
	.I2(r_4[0]),
	.I3(r_4[1]),
	.O(un26_r_lt0)
);
defparam un26_r_lt0_cZ.INIT=16'h08AE;
// @7:143
  MUXCY_L \b18_cry_cZ[28]  (
	.DI(b18_lt28),
	.CI(b18_cry[26]),
	.S(b18_df28),
	.LO(b18_cry[28])
);
// @7:143
  MUXCY_L \b18_cry_cZ[26]  (
	.DI(b18_lt26),
	.CI(b18_cry[24]),
	.S(b18_df26),
	.LO(b18_cry[26])
);
// @7:143
  MUXCY_L \b18_cry_cZ[24]  (
	.DI(b18_lt24),
	.CI(b18_cry[22]),
	.S(b18_df24),
	.LO(b18_cry[24])
);
// @7:143
  MUXCY_L \b18_cry_cZ[22]  (
	.DI(b18_lt22),
	.CI(b18_cry[20]),
	.S(b18_df22),
	.LO(b18_cry[22])
);
// @7:143
  MUXCY_L \b18_cry_cZ[20]  (
	.DI(b18_lt20),
	.CI(b18_cry[18]),
	.S(b18_df20),
	.LO(b18_cry[20])
);
// @7:143
  MUXCY_L \b18_cry_cZ[18]  (
	.DI(b18_lt18),
	.CI(b18_cry[16]),
	.S(b18_df18),
	.LO(b18_cry[18])
);
// @7:143
  LUT4 b18_lt18_cZ (
	.I0(m_2[19]),
	.I1(m_2[18]),
	.I2(r_4[19]),
	.I3(r_4[18]),
	.O(b18_lt18)
);
defparam b18_lt18_cZ.INIT=16'h7150;
// @7:143
  MUXCY_L \b18_cry_cZ[16]  (
	.DI(b18_lt16),
	.CI(b18_cry[14]),
	.S(b18_df16),
	.LO(b18_cry[16])
);
// @7:143
  LUT4 b18_lt16_cZ (
	.I0(m_2[16]),
	.I1(m_2[17]),
	.I2(r_4[16]),
	.I3(r_4[17]),
	.O(b18_lt16)
);
defparam b18_lt16_cZ.INIT=16'h7310;
// @7:143
  MUXCY_L \b18_cry_cZ[14]  (
	.DI(b18_lt14),
	.CI(b18_cry[12]),
	.S(b18_df14),
	.LO(b18_cry[14])
);
// @7:143
  LUT4 b18_lt14_cZ (
	.I0(m_2[14]),
	.I1(m_2[15]),
	.I2(r_4[14]),
	.I3(r_4[15]),
	.O(b18_lt14)
);
defparam b18_lt14_cZ.INIT=16'h7310;
// @7:143
  MUXCY_L \b18_cry_cZ[12]  (
	.DI(b18_lt12),
	.CI(b18_cry[10]),
	.S(b18_df12),
	.LO(b18_cry[12])
);
// @7:143
  LUT4 b18_lt12_cZ (
	.I0(m_2[12]),
	.I1(m_2[13]),
	.I2(r_4[12]),
	.I3(r_4[13]),
	.O(b18_lt12)
);
defparam b18_lt12_cZ.INIT=16'h7310;
// @7:143
  MUXCY_L \b18_cry_cZ[10]  (
	.DI(b18_lt10),
	.CI(b18_cry[8]),
	.S(b18_df10),
	.LO(b18_cry[10])
);
// @7:143
  LUT4 b18_lt10_cZ (
	.I0(m_2[10]),
	.I1(m_2[11]),
	.I2(r_4[11]),
	.I3(r_4[10]),
	.O(b18_lt10)
);
defparam b18_lt10_cZ.INIT=16'h7130;
// @7:143
  MUXCY_L \b18_cry_cZ[8]  (
	.DI(b18_lt8),
	.CI(b18_cry[6]),
	.S(b18_df8),
	.LO(b18_cry[8])
);
// @7:143
  LUT4 b18_lt8_cZ (
	.I0(m_2[8]),
	.I1(m_2[9]),
	.I2(r_4[8]),
	.I3(r_4[9]),
	.O(b18_lt8)
);
defparam b18_lt8_cZ.INIT=16'h7310;
// @7:143
  MUXCY_L \b18_cry_cZ[6]  (
	.DI(b18_lt6),
	.CI(b18_cry[4]),
	.S(b18_df6),
	.LO(b18_cry[6])
);
// @7:143
  LUT4 b18_lt6_cZ (
	.I0(m_2[7]),
	.I1(m_2[6]),
	.I2(r_4[6]),
	.I3(r_4[7]),
	.O(b18_lt6)
);
defparam b18_lt6_cZ.INIT=16'h7510;
// @7:143
  MUXCY_L \b18_cry_cZ[4]  (
	.DI(b18_lt4),
	.CI(b18_cry[2]),
	.S(b18_df4),
	.LO(b18_cry[4])
);
// @7:143
  LUT4 b18_lt4_cZ (
	.I0(m_2[4]),
	.I1(m_2[5]),
	.I2(r_4[4]),
	.I3(r_4[5]),
	.O(b18_lt4)
);
defparam b18_lt4_cZ.INIT=16'h7310;
// @7:143
  MUXCY_L \b18_cry_cZ[2]  (
	.DI(b18_lt2),
	.CI(b18_cry[0]),
	.S(b18_df2),
	.LO(b18_cry[2])
);
// @7:143
  LUT4 b18_lt2_cZ (
	.I0(m_2[2]),
	.I1(m_2[3]),
	.I2(r_4[3]),
	.I3(N_28),
	.O(b18_lt2)
);
defparam b18_lt2_cZ.INIT=16'h7130;
// @7:143
  MUXCY_L \b18_cry_cZ[0]  (
	.DI(b18_lt0),
	.CI(GND),
	.S(b18_df0),
	.LO(b18_cry[0])
);
// @7:143
  LUT4 b18_lt0_cZ (
	.I0(m_2[1]),
	.I1(m_2[0]),
	.I2(r_4[0]),
	.I3(r_4[1]),
	.O(b18_lt0)
);
defparam b18_lt0_cZ.INIT=16'h7510;
// @7:118
  MUXCY_L \un11_r_cry_cZ[28]  (
	.DI(un11_r_lt28),
	.CI(un11_r_cry[26]),
	.S(un11_r_df28),
	.LO(un11_r_cry[28])
);
// @7:118
  MUXCY_L \un11_r_cry_cZ[26]  (
	.DI(un11_r_lt26),
	.CI(un11_r_cry[24]),
	.S(un11_r_df26),
	.LO(un11_r_cry[26])
);
// @7:118
  MUXCY_L \un11_r_cry_cZ[24]  (
	.DI(un11_r_lt24),
	.CI(un11_r_cry[22]),
	.S(un11_r_df24),
	.LO(un11_r_cry[24])
);
// @7:118
  MUXCY_L \un11_r_cry_cZ[22]  (
	.DI(un11_r_lt22),
	.CI(un11_r_cry[20]),
	.S(un11_r_df22),
	.LO(un11_r_cry[22])
);
// @7:118
  MUXCY_L \un11_r_cry_cZ[20]  (
	.DI(un11_r_lt20),
	.CI(un11_r_cry[18]),
	.S(un11_r_df20),
	.LO(un11_r_cry[20])
);
// @7:118
  MUXCY_L \un11_r_cry_cZ[18]  (
	.DI(un11_r_lt18),
	.CI(un11_r_cry[16]),
	.S(un11_r_df18),
	.LO(un11_r_cry[18])
);
// @7:118
  LUT4 un11_r_lt18_cZ (
	.I0(m_2[19]),
	.I1(m_2[18]),
	.I2(r_4[19]),
	.I3(r_4[18]),
	.O(un11_r_lt18)
);
defparam un11_r_lt18_cZ.INIT=16'h0A8E;
// @7:118
  MUXCY_L \un11_r_cry_cZ[16]  (
	.DI(un11_r_lt16),
	.CI(un11_r_cry[14]),
	.S(un11_r_df16),
	.LO(un11_r_cry[16])
);
// @7:118
  LUT4 un11_r_lt16_cZ (
	.I0(m_2[16]),
	.I1(m_2[17]),
	.I2(r_4[16]),
	.I3(r_4[17]),
	.O(un11_r_lt16)
);
defparam un11_r_lt16_cZ.INIT=16'h08CE;
// @7:118
  MUXCY_L \un11_r_cry_cZ[14]  (
	.DI(un11_r_lt14),
	.CI(un11_r_cry[12]),
	.S(un11_r_df14),
	.LO(un11_r_cry[14])
);
// @7:118
  LUT4 un11_r_lt14_cZ (
	.I0(m_2[14]),
	.I1(m_2[15]),
	.I2(r_4[14]),
	.I3(r_4[15]),
	.O(un11_r_lt14)
);
defparam un11_r_lt14_cZ.INIT=16'h08CE;
// @7:118
  MUXCY_L \un11_r_cry_cZ[12]  (
	.DI(un11_r_lt12),
	.CI(un11_r_cry[10]),
	.S(un11_r_df12),
	.LO(un11_r_cry[12])
);
// @7:118
  LUT4 un11_r_lt12_cZ (
	.I0(m_2[12]),
	.I1(m_2[13]),
	.I2(r_4[12]),
	.I3(r_4[13]),
	.O(un11_r_lt12)
);
defparam un11_r_lt12_cZ.INIT=16'h08CE;
// @7:118
  MUXCY_L \un11_r_cry_cZ[10]  (
	.DI(un11_r_lt10),
	.CI(un11_r_cry[8]),
	.S(un11_r_df10),
	.LO(un11_r_cry[10])
);
// @7:118
  LUT4 un11_r_lt10_cZ (
	.I0(m_2[10]),
	.I1(m_2[11]),
	.I2(r_4[11]),
	.I3(r_4[10]),
	.O(un11_r_lt10)
);
defparam un11_r_lt10_cZ.INIT=16'h0C8E;
// @7:118
  MUXCY_L \un11_r_cry_cZ[8]  (
	.DI(un11_r_lt8),
	.CI(un11_r_cry[6]),
	.S(un11_r_df8),
	.LO(un11_r_cry[8])
);
// @7:118
  LUT4 un11_r_lt8_cZ (
	.I0(m_2[8]),
	.I1(m_2[9]),
	.I2(r_4[8]),
	.I3(r_4[9]),
	.O(un11_r_lt8)
);
defparam un11_r_lt8_cZ.INIT=16'h08CE;
// @7:118
  MUXCY_L \un11_r_cry_cZ[6]  (
	.DI(un11_r_lt6),
	.CI(un11_r_cry[4]),
	.S(un11_r_df6),
	.LO(un11_r_cry[6])
);
// @7:118
  LUT4 un11_r_lt6_cZ (
	.I0(m_2[7]),
	.I1(m_2[6]),
	.I2(r_4[6]),
	.I3(r_4[7]),
	.O(un11_r_lt6)
);
defparam un11_r_lt6_cZ.INIT=16'h08AE;
// @7:118
  MUXCY_L \un11_r_cry_cZ[4]  (
	.DI(un11_r_lt4),
	.CI(un11_r_cry[2]),
	.S(un11_r_df4),
	.LO(un11_r_cry[4])
);
// @7:118
  LUT4 un11_r_lt4_cZ (
	.I0(m_2[4]),
	.I1(m_2[5]),
	.I2(r_4[4]),
	.I3(r_4[5]),
	.O(un11_r_lt4)
);
defparam un11_r_lt4_cZ.INIT=16'h08CE;
// @7:118
  MUXCY_L \un11_r_cry_cZ[2]  (
	.DI(un11_r_lt2),
	.CI(un11_r_cry[0]),
	.S(un11_r_df2),
	.LO(un11_r_cry[2])
);
// @7:118
  LUT4 un11_r_lt2_cZ (
	.I0(m_2[2]),
	.I1(m_2[3]),
	.I2(r_4[3]),
	.I3(N_28),
	.O(un11_r_lt2)
);
defparam un11_r_lt2_cZ.INIT=16'h0C8E;
// @7:118
  MUXCY_L \un11_r_cry_cZ[0]  (
	.DI(un11_r_lt0),
	.CI(GND),
	.S(un11_r_df0),
	.LO(un11_r_cry[0])
);
// @7:118
  LUT4 un11_r_lt0_cZ (
	.I0(m_2[1]),
	.I1(m_2[0]),
	.I2(r_4[0]),
	.I3(r_4[1]),
	.O(un11_r_lt0)
);
defparam un11_r_lt0_cZ.INIT=16'h08AE;
// @7:128
  MUXCY_L un14_r_0_I_75 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[3]),
	.S(un14_r_0_N_7),
	.LO(un14_r_0_data_tmp[4])
);
// @7:128
  MUXCY_L un14_r_0_I_67 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[0]),
	.S(un14_r_0_N_14),
	.LO(un14_r_0_data_tmp[1])
);
// @7:128
  MUXCY_L un14_r_0_I_59 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[1]),
	.S(un14_r_0_N_21),
	.LO(un14_r_0_data_tmp[2])
);
// @7:128
  MUXCY_L un14_r_0_I_51 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[2]),
	.S(un14_r_0_N_28),
	.LO(un14_r_0_data_tmp[3])
);
// @7:128
  MUXCY_L un14_r_0_I_43 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[7]),
	.S(un14_r_0_N_35),
	.LO(un14_r_0_data_tmp[8])
);
// @7:128
  MUXCY_L un14_r_0_I_35 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[4]),
	.S(un14_r_0_N_42),
	.LO(un14_r_0_data_tmp[5])
);
// @7:128
  MUXCY_L un14_r_0_I_27 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[5]),
	.S(un14_r_0_N_49),
	.LO(un14_r_0_data_tmp[6])
);
// @7:128
  MUXCY_L un14_r_0_I_19 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[6]),
	.S(un14_r_0_N_56),
	.LO(un14_r_0_data_tmp[7])
);
// @7:128
  MUXCY_L un14_r_0_I_11 (
	.DI(GND),
	.CI(un14_r_0_data_tmp[8]),
	.S(un14_r_0_N_63),
	.LO(un14_r_0_data_tmp[9])
);
// @7:128
  MUXCY_L un14_r_0_I_1 (
	.DI(GND),
	.CI(VCC),
	.S(un14_r_0_N_70),
	.LO(un14_r_0_data_tmp[0])
);
// @7:47
  LUT4 \d_cnst_sn.reg0_28_5_2426_a6_1_1_lut6_2_o6  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(reg3_1_1[21]),
	.O(\d_cnst_sn.reg0_28_5_2426_a6_1_1 )
);
defparam \d_cnst_sn.reg0_28_5_2426_a6_1_1_lut6_2_o6 .INIT=16'h0100;
// @7:47
  LUT3 \d_cnst_sn.reg0_28_5_2426_a6_1_1_lut6_2_o5  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.O(\d_cnst_sn.reg0_28_12_2195_a6_1_2_0 )
);
defparam \d_cnst_sn.reg0_28_5_2426_a6_1_1_lut6_2_o5 .INIT=8'h01;
// @7:47
  LUT4 \d_cnst_sn.reg0_28_9_2294_a6_1_1_lut6_2_o6  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(reg3_1_1[25]),
	.O(\d_cnst_sn.reg0_28_9_2294_a6_1_1 )
);
defparam \d_cnst_sn.reg0_28_9_2294_a6_1_1_lut6_2_o6 .INIT=16'h0100;
// @7:47
  LUT4 \d_cnst_sn.reg0_28_9_2294_a6_1_1_lut6_2_o5  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(reg3_1_1[26]),
	.O(\d_cnst_sn.reg0_28_10_2261_a6_1_1 )
);
defparam \d_cnst_sn.reg0_28_9_2294_a6_1_1_lut6_2_o5 .INIT=16'h0100;
// @7:97
  LUT2 \d_cnst_sn.r_4_2_a1_lut6_2_o6[3]  (
	.I0(reg1[3]),
	.I1(inf_abs0_2[30]),
	.O(r_4_2_a1_lut6_2_O6[3])
);
defparam \d_cnst_sn.r_4_2_a1_lut6_2_o6[3] .INIT=4'h1;
// @7:97
  LUT2 \d_cnst_sn.r_4_2_a1_lut6_2_o5[3]  (
	.I0(reg1[4]),
	.I1(inf_abs0_2[30]),
	.O(r_4_2_a1_lut6_2_O5[3])
);
defparam \d_cnst_sn.r_4_2_a1_lut6_2_o5[3] .INIT=4'h1;
// @7:47
  LUT4 \d_cnst_sn.reg0_28_7_2360_a6_1_1_lut6_2_o6  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(reg3_1_1[23]),
	.O(\d_cnst_sn.reg0_28_7_2360_a6_1_1 )
);
defparam \d_cnst_sn.reg0_28_7_2360_a6_1_1_lut6_2_o6 .INIT=16'h0100;
// @7:47
  LUT2 \d_cnst_sn.reg0_28_7_2360_a6_1_1_lut6_2_o5  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.O(N_3873_2)
);
defparam \d_cnst_sn.reg0_28_7_2360_a6_1_1_lut6_2_o5 .INIT=4'h1;
  LUT2 \d_cnst_sn.g0_0_0_a5_0_0_lut6_2_o6  (
	.I0(datai[31]),
	.I1(inf_abs0_2[20]),
	.O(\d_cnst_sn.g0_0_0_a5_0_0 )
);
defparam \d_cnst_sn.g0_0_0_a5_0_0_lut6_2_o6 .INIT=4'h8;
  LUT3 \d_cnst_sn.g0_0_0_a5_0_0_lut6_2_o5  (
	.I0(datai[20]),
	.I1(state[0]),
	.I2(inf_abs0_2[20]),
	.O(ir_3[20])
);
defparam \d_cnst_sn.g0_0_0_a5_0_0_lut6_2_o5 .INIT=8'hE2;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_1052_i_a6_2_0_lut6_2_o6  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.I2(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 )
);
defparam \d_cnst_sn.addr_20_iv_1052_i_a6_2_0_lut6_2_o6 .INIT=8'h80;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_1052_i_a6_2_0_lut6_2_o5  (
	.I0(datai[30]),
	.I1(state[0]),
	.I2(inf_abs0_2[30]),
	.O(ir_3[30])
);
defparam \d_cnst_sn.addr_20_iv_1052_i_a6_2_0_lut6_2_o5 .INIT=8'hE2;
// @7:47
  LUT2 \d_cnst_sn.addr_20_iv_1052_i_a6_1_0_lut6_2_o6  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.O(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 )
);
defparam \d_cnst_sn.addr_20_iv_1052_i_a6_1_0_lut6_2_o6 .INIT=4'h2;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_1052_i_a6_1_0_lut6_2_o5  (
	.I0(datai[31]),
	.I1(state[0]),
	.I2(inf_abs0_2[31]),
	.O(ir_3[31])
);
defparam \d_cnst_sn.addr_20_iv_1052_i_a6_1_0_lut6_2_o5 .INIT=8'hE2;
// @7:47
  LUT3 \d_cnst_sn.reg0_28_10_2261_a6_1_0_lut6_2_o6  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.O(\d_cnst_sn.reg0_28_2526_a5_1_0 )
);
defparam \d_cnst_sn.reg0_28_10_2261_a6_1_0_lut6_2_o6 .INIT=8'h01;
// @7:47
  LUT4 \d_cnst_sn.reg0_28_10_2261_a6_1_0_lut6_2_o5  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.g0_0_0_a5_2 )
);
defparam \d_cnst_sn.reg0_28_10_2261_a6_1_0_lut6_2_o5 .INIT=16'h0008;
// @7:47
  LUT4 \d_cnst_sn.g0_2_lut6_2_o6  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg0_N_13_0 )
);
defparam \d_cnst_sn.g0_2_lut6_2_o6 .INIT=16'h003E;
// @7:47
  LUT3 \d_cnst_sn.g0_2_lut6_2_o5  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg0_m8_e_0 )
);
defparam \d_cnst_sn.g0_2_lut6_2_o5 .INIT=8'h07;
// @7:47
  LUT4 \d_cnst_sn.reg0_28_8_2327_a6_1_1_lut6_2_o6  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(reg3_1_1[24]),
	.O(\d_cnst_sn.reg0_28_8_2327_a6_1_1 )
);
defparam \d_cnst_sn.reg0_28_8_2327_a6_1_1_lut6_2_o6 .INIT=16'h0100;
// @7:47
  LUT3 \d_cnst_sn.reg0_28_8_2327_a6_1_1_lut6_2_o5  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg1_16_8_1837_2_tz )
);
defparam \d_cnst_sn.reg0_28_8_2327_a6_1_1_lut6_2_o5 .INIT=8'hF8;
// @7:86
  LUT2 \d_cnst_sn.r_4_2_RNIBJSG2_o6[18]  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[28]),
	.O(N_527_i)
);
defparam \d_cnst_sn.r_4_2_RNIBJSG2_o6[18] .INIT=4'h4;
// @7:86
  LUT5 \d_cnst_sn.r_4_2_RNIBJSG2_o5[18]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[18]),
	.I4(reg3_1_1[19]),
	.O(\d_cnst_sn.reg0_28_0 [19])
);
defparam \d_cnst_sn.r_4_2_RNIBJSG2_o5[18] .INIT=32'hFFDF2202;
// @7:47
  LUT4 \d_cnst_sn.addr_20_iv_6_863_i_0_lut6_2_o6  (
	.I0(reg3[19]),
	.I1(state[0]),
	.I2(inf_abs0_2[19]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_6_863_i_0 )
);
defparam \d_cnst_sn.addr_20_iv_6_863_i_0_lut6_2_o6 .INIT=16'h111D;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_6_863_i_0_lut6_2_o5  (
	.I0(datai[28]),
	.I1(state[0]),
	.I2(inf_abs0_2[28]),
	.O(ir_3[28])
);
defparam \d_cnst_sn.addr_20_iv_6_863_i_0_lut6_2_o5 .INIT=8'hE2;
// @7:106
  LUT2 \d_cnst_sn.g0_2_0_i2_lut6_2_o6  (
	.I0(inf_abs0_2[27]),
	.I1(inf_abs0_2[28]),
	.O(g0_2_0_i2_lut6_2_O6)
);
defparam \d_cnst_sn.g0_2_0_i2_lut6_2_o6 .INIT=4'h1;
// @7:106
  LUT4 \d_cnst_sn.g0_2_0_i2_lut6_2_o5  (
	.I0(reg3[18]),
	.I1(state[0]),
	.I2(inf_abs0_2[18]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_5_890_i_0 )
);
defparam \d_cnst_sn.g0_2_0_i2_lut6_2_o5 .INIT=16'h111D;
// @7:47
  LUT4 \d_cnst_sn.addr_20_iv_4_917_i_0_lut6_2_o6  (
	.I0(reg3[17]),
	.I1(state[0]),
	.I2(inf_abs0_2[17]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_4_917_i_0 )
);
defparam \d_cnst_sn.addr_20_iv_4_917_i_0_lut6_2_o6 .INIT=16'h111D;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_4_917_i_0_lut6_2_o5  (
	.I0(datai[17]),
	.I1(state[0]),
	.I2(inf_abs0_2[17]),
	.O(ir_3[17])
);
defparam \d_cnst_sn.addr_20_iv_4_917_i_0_lut6_2_o5 .INIT=8'hE2;
// @7:47
  LUT2 \d_cnst_sn.g0_3_o2_lut6_2_o6  (
	.I0(inf_abs0_2[27]),
	.I1(inf_abs0_2[28]),
	.O(N_7)
);
defparam \d_cnst_sn.g0_3_o2_lut6_2_o6 .INIT=4'hE;
// @7:47
  LUT4 \d_cnst_sn.g0_3_o2_lut6_2_o5  (
	.I0(reg3[16]),
	.I1(state[0]),
	.I2(inf_abs0_2[16]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_3_944_i_0 )
);
defparam \d_cnst_sn.g0_3_o2_lut6_2_o5 .INIT=16'h111D;
// @7:47
  LUT4 \d_cnst_sn.addr_20_iv_0_1025_i_0_lut6_2_o6  (
	.I0(reg3[13]),
	.I1(state[0]),
	.I2(inf_abs0_2[13]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_0_1025_i_0 )
);
defparam \d_cnst_sn.addr_20_iv_0_1025_i_0_lut6_2_o6 .INIT=16'h111D;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_0_1025_i_0_lut6_2_o5  (
	.I0(datai[13]),
	.I1(state[0]),
	.I2(inf_abs0_2[13]),
	.O(ir_3[13])
);
defparam \d_cnst_sn.addr_20_iv_0_1025_i_0_lut6_2_o5 .INIT=8'hE2;
// @7:47
  LUT4 \d_cnst_sn.addr_20_iv_1052_i_0_lut6_2_o6  (
	.I0(reg3[12]),
	.I1(state[0]),
	.I2(inf_abs0_2[12]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_1052_i_0 )
);
defparam \d_cnst_sn.addr_20_iv_1052_i_0_lut6_2_o6 .INIT=16'h111D;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_1052_i_0_lut6_2_o5  (
	.I0(datai[12]),
	.I1(state[0]),
	.I2(inf_abs0_2[12]),
	.O(ir_3[12])
);
defparam \d_cnst_sn.addr_20_iv_1052_i_0_lut6_2_o5 .INIT=8'hE2;
// @7:47
  LUT4 \d_cnst_sn.addr_20_iv_1_998_i_0_lut6_2_o6  (
	.I0(reg3[14]),
	.I1(state[0]),
	.I2(inf_abs0_2[14]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_1_998_i_0 )
);
defparam \d_cnst_sn.addr_20_iv_1_998_i_0_lut6_2_o6 .INIT=16'h111D;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_1_998_i_0_lut6_2_o5  (
	.I0(datai[14]),
	.I1(state[0]),
	.I2(inf_abs0_2[14]),
	.O(ir_3[14])
);
defparam \d_cnst_sn.addr_20_iv_1_998_i_0_lut6_2_o5 .INIT=8'hE2;
// @7:47
  LUT4 \d_cnst_sn.addr_20_iv_2_971_i_0_lut6_2_o6  (
	.I0(reg3[15]),
	.I1(state[0]),
	.I2(inf_abs0_2[15]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.addr_20_iv_2_971_i_0 )
);
defparam \d_cnst_sn.addr_20_iv_2_971_i_0_lut6_2_o6 .INIT=16'h111D;
// @7:47
  LUT3 \d_cnst_sn.addr_20_iv_2_971_i_0_lut6_2_o5  (
	.I0(datai[15]),
	.I1(state[0]),
	.I2(inf_abs0_2[15]),
	.O(ir_3[15])
);
defparam \d_cnst_sn.addr_20_iv_2_971_i_0_lut6_2_o5 .INIT=8'hE2;
// @7:47
  LUT4 \d_cnst_sn.reg0_28_6_2393_a6_1_1_lut6_2_o6  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(reg3_1_1[22]),
	.O(\d_cnst_sn.reg0_28_6_2393_a6_1_1 )
);
defparam \d_cnst_sn.reg0_28_6_2393_a6_1_1_lut6_2_o6 .INIT=16'h0100;
// @7:47
  LUT3 \d_cnst_sn.reg0_28_6_2393_a6_1_1_lut6_2_o5  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.O(\d_cnst_sn.b60_0 )
);
defparam \d_cnst_sn.reg0_28_6_2393_a6_1_1_lut6_2_o5 .INIT=8'h02;
// @7:47
  LUT2 \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_o6  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[31]),
	.O(N_512_i)
);
defparam \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_o6 .INIT=4'h2;
// @7:47
  LUT3 \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_o5  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg0_m9_i_a3_0 )
);
defparam \d_cnst_sn.reg0_28_10_2261_a6_3_2_lut6_2_o5 .INIT=8'h06;
// @7:74
  LUT5 \d_cnst_sn.reg0_28_0_lut6_2_o6[20]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.I3(r_4[19]),
	.I4(reg3_1_1[20]),
	.O(\d_cnst_sn.reg0_28_0 [20])
);
defparam \d_cnst_sn.reg0_28_0_lut6_2_o6[20] .INIT=32'hFFDF2202;
// @7:74
  LUT3 \d_cnst_sn.reg0_28_0_lut6_2_o5[20]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[28]),
	.O(\d_cnst_sn.reg0_28_7_a0_0 [9])
);
defparam \d_cnst_sn.reg0_28_0_lut6_2_o5[20] .INIT=8'h02;
// @7:74
  LUT3 \d_cnst_sn.reg0_28_a2_0_lut6_2_o6[2]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg1_16_a2_0 [5])
);
defparam \d_cnst_sn.reg0_28_a2_0_lut6_2_o6[2] .INIT=8'hF1;
// @7:74
  LUT2 \d_cnst_sn.reg0_28_a2_0_lut6_2_o5[2]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[31]),
	.O(N_3913)
);
defparam \d_cnst_sn.reg0_28_a2_0_lut6_2_o5[2] .INIT=4'hD;
// @7:74
  LUT3 \d_cnst_sn.reg2_16_11_a0_0_lut6_2_o6[31]  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg2_N_3_mux )
);
defparam \d_cnst_sn.reg2_16_11_a0_0_lut6_2_o6[31] .INIT=8'hF1;
// @7:74
  LUT5 \d_cnst_sn.reg2_16_11_a0_0_lut6_2_o5[31]  (
	.I0(reg3[0]),
	.I1(inf_abs0_2[19]),
	.I2(inf_abs0_2[20]),
	.I3(inf_abs0_2[31]),
	.I4(m_2[0]),
	.O(N_1335)
);
defparam \d_cnst_sn.reg2_16_11_a0_0_lut6_2_o5[31] .INIT=32'hFFFB0008;
// @7:179
  LUT3 \d_cnst_sn.b64_0_lut6_2_o6  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.O(\d_cnst_sn.b64_0 )
);
defparam \d_cnst_sn.b64_0_lut6_2_o6 .INIT=8'h04;
// @7:179
  LUT2 \d_cnst_sn.b64_0_lut6_2_o5  (
	.I0(inf_abs0_2[31]),
	.I1(inf_abs0_2[27]),
	.O(N_526_i)
);
defparam \d_cnst_sn.b64_0_lut6_2_o5 .INIT=4'h4;
// @7:105
  LUT4 \d_cnst_sn.m_2_lut6_2_o6[30]  (
	.I0(datai[30]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[30])
);
defparam \d_cnst_sn.m_2_lut6_2_o6[30] .INIT=16'h2220;
// @7:105
  LUT4 \d_cnst_sn.m_2_lut6_2_o5[30]  (
	.I0(datai[31]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2[31])
);
defparam \d_cnst_sn.m_2_lut6_2_o5[30] .INIT=16'h2220;
// @7:184
  LUT3 \d_cnst_sn.reg0_28_sn_m6_lut6_2_o6  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.O(N_3916)
);
defparam \d_cnst_sn.reg0_28_sn_m6_lut6_2_o6 .INIT=8'h06;
// @7:184
  LUT3 \d_cnst_sn.reg0_28_sn_m6_lut6_2_o5  (
	.I0(b),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.O(reg0_28_sn_m6_lut6_2_O5)
);
defparam \d_cnst_sn.reg0_28_sn_m6_lut6_2_o5 .INIT=8'h20;
// @7:47
  LUT4 \d_cnst_sn.reg0_m9_i_a0_0_lut6_2_o6  (
	.I0(b),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[27]),
	.O(\d_cnst_sn.reg0_m9_i_a0_0 )
);
defparam \d_cnst_sn.reg0_m9_i_a0_0_lut6_2_o6 .INIT=16'h040C;
// @7:47
  LUT2 \d_cnst_sn.reg0_m9_i_a0_0_lut6_2_o5  (
	.I0(state[0]),
	.I1(inf_abs0_2[27]),
	.O(N_2660_2)
);
defparam \d_cnst_sn.reg0_m9_i_a0_0_lut6_2_o5 .INIT=4'h8;
// @7:74
  LUT4 \d_cnst_sn.reg0_28_a1_1_lut6_2_o6[7]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.O(N_3910)
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_o6[7] .INIT=16'h0002;
// @7:74
  LUT4 \d_cnst_sn.reg0_28_a1_1_lut6_2_o5[7]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.g0_3_a2_2 )
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_o5[7] .INIT=16'h0008;
// @7:74
  LUT4 \d_cnst_sn.reg0_28_a1_1_lut6_2_o6[2]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.reg0_28_a1_1 [4])
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_o6[2] .INIT=16'h0800;
// @7:74
  LUT4 \d_cnst_sn.reg0_28_a1_1_lut6_2_o5[2]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg0_28_9_2294_a6_3_0 )
);
defparam \d_cnst_sn.reg0_28_a1_1_lut6_2_o5[2] .INIT=16'h0002;
// @7:74
  LUT4 \d_cnst_sn.reg0_28_a0_1_lut6_2_o6[7]  (
	.I0(inf_abs0_2[20]),
	.I1(inf_abs0_2[21]),
	.I2(inf_abs0_2[22]),
	.I3(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg0_28_a0_1 [7])
);
defparam \d_cnst_sn.reg0_28_a0_1_lut6_2_o6[7] .INIT=16'hFF01;
// @7:74
  LUT4 \d_cnst_sn.reg0_28_a0_1_lut6_2_o5[7]  (
	.I0(inf_abs0_2[21]),
	.I1(inf_abs0_2[22]),
	.I2(inf_abs0_2[31]),
	.I3(inf_abs0_2[28]),
	.O(\d_cnst_sn.reg1_16_a0_1 [3])
);
defparam \d_cnst_sn.reg0_28_a0_1_lut6_2_o5[7] .INIT=16'h0008;
// @7:243
  LUT4 \d_cnst_sn.m_2_i_lut6_2_o6[31]  (
	.I0(datai[31]),
	.I1(inf_abs0_2[31]),
	.I2(inf_abs0_2[27]),
	.I3(inf_abs0_2[28]),
	.O(m_2_i[31])
);
defparam \d_cnst_sn.m_2_i_lut6_2_o6[31] .INIT=16'hDDDF;
// @7:243
  LUT3 \d_cnst_sn.m_2_i_lut6_2_o5[31]  (
	.I0(datai[31]),
	.I1(state[0]),
	.I2(inf_abs0_2[31]),
	.O(ir_3_fast[31])
);
defparam \d_cnst_sn.m_2_i_lut6_2_o5[31] .INIT=8'hE2;
// @7:184
  LUT4 \d_cnst_sn.reg0_28_sn_m4_lut6_2_o6  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[31]),
	.O(N_1033)
);
defparam \d_cnst_sn.reg0_28_sn_m4_lut6_2_o6 .INIT=16'hFF35;
// @7:184
  LUT5 \d_cnst_sn.reg0_28_sn_m4_lut6_2_o5  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg2_16_11_1_tz [28])
);
defparam \d_cnst_sn.reg0_28_sn_m4_lut6_2_o5 .INIT=32'hFFFFFACF;
// @7:74
  LUT5 \d_cnst_sn.un1_state_1_1_a6_0_lut6_2_o6  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.O(N_1892)
);
defparam \d_cnst_sn.un1_state_1_1_a6_0_lut6_2_o6 .INIT=32'h0000E000;
// @7:74
  LUT5 \d_cnst_sn.un1_state_1_1_a6_0_lut6_2_o5  (
	.I0(inf_abs0_2[19]),
	.I1(inf_abs0_2[20]),
	.I2(inf_abs0_2[21]),
	.I3(inf_abs0_2[22]),
	.I4(inf_abs0_2[31]),
	.O(\d_cnst_sn.reg2_16_0_1_tz [28])
);
defparam \d_cnst_sn.un1_state_1_1_a6_0_lut6_2_o5 .INIT=32'hFFFFF53F;
// @7:143
  LUT4 b18_df30_lut6_2_o6 (
	.I0(m_2_i[31]),
	.I1(r_4[30]),
	.I2(m_2[30]),
	.I3(r_4_i[31]),
	.O(b18_df30)
);
defparam b18_df30_lut6_2_o6.INIT=16'h8241;
// @7:143
  LUT4 b18_df30_lut6_2_o5 (
	.I0(m_2_i[31]),
	.I1(r_4[30]),
	.I2(m_2[30]),
	.I3(r_4_i[31]),
	.O(b18_lt30)
);
defparam b18_df30_lut6_2_o5.INIT=16'h5D04;
// @7:118
  LUT4 un11_r_df30_lut6_2_o6 (
	.I0(m_2_i[31]),
	.I1(r_4[30]),
	.I2(m_2[30]),
	.I3(r_4_i[31]),
	.O(un11_r_df30)
);
defparam un11_r_df30_lut6_2_o6.INIT=16'h8241;
// @7:118
  LUT4 un11_r_df30_lut6_2_o5 (
	.I0(m_2_i[31]),
	.I1(r_4[30]),
	.I2(m_2[30]),
	.I3(r_4_i[31]),
	.O(un11_r_lt30)
);
defparam un11_r_df30_lut6_2_o5.INIT=16'h20BA;
endmodule