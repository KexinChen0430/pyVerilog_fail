module t (/*AUTOARG*/
   // Inputs
   clk
   );
   input clk;
   reg [pkg11::PARAM1 : 0] bus11;
   reg [pkg11::PARAM2 : 0] bus12;
   reg [pkg11::PARAM3 : 0] bus13;
   reg [pkg21::PARAM1 : 0] bus21;
   reg [pkg21::PARAM2 : 0] bus22;
   reg [pkg21::PARAM3 : 0] bus23;
   reg [pkg31::PARAM1 : 0] bus31;
   reg [pkg31::PARAM2 : 0] bus32;
   reg [pkg31::PARAM3 : 0] bus33;
   initial begin
      $write("*-* All Finished *-*\n");
      $finish;
   end
endmodule