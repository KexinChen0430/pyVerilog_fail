module INBUF (
	(* iopad_external_pin *)
	input PAD,
	output Y
);
	assign Y = PAD;
endmodule