module my_NDI1MUX_NDI1 (input clk, input [31:0] din, output [7:0] dout);
    parameter LOC = "SLICE_X6Y100";
    wire [3:0] q31;
    (* LOC=LOC, BEL="D6LUT" *)
    SRLC32E #(
            .INIT(32'h00000000),
            .IS_CLK_INVERTED(1'b0)
        ) lutd (
            .Q(dout[0]),
            .Q31(q31[3]),
            .A(din[4:0]),
            .CE(din[5]),
            .CLK(din[6]),
            .D(din[7]));
    (* LOC=LOC, BEL="C6LUT" *)
    SRLC32E #(
            .INIT(32'h00000000),
            .IS_CLK_INVERTED(1'b0)
        ) lutc (
            .Q(dout[1]),
            .Q31(q31[2]),
            .A(din[12:8]),
            .CE(din[5]),
            .CLK(din[6]),
            .D(din[15]));
    (* LOC=LOC, BEL="B6LUT" *)
    SRLC32E #(
            .INIT(32'h00000000),
            .IS_CLK_INVERTED(1'b0)
        ) lutb (
            .Q(dout[2]),
            .Q31(q31[1]),
            .A(din[20:16]),
            .CE(din[5]),
            .CLK(din[6]),
            //.D(din[23]));
            .D(q31[2]));
    (* LOC=LOC, BEL="A6LUT" *)
    SRLC32E #(
            .INIT(32'h00000000),
            .IS_CLK_INVERTED(1'b0)
        ) luta (
            .Q(dout[3]),
            .Q31(q31[0]),
            .A(din[28:24]),
            .CE(din[5]),
            .CLK(din[6]),
            //.D(din[31]));
            .D(q31[2]));
endmodule