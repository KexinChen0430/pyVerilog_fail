module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_eda
		inst_eda_e inst_eda (
		);
		// End of Generated Instance Port Map for inst_eda
		// Generated Instance Port Map for inst_edb
		inst_edb_e inst_edb (
		);
		// End of Generated Instance Port Map for inst_edb
endmodule