module OB(input I,
	(* iopad_external_pin *) output O);
	assign O = I;
endmodule