module adder (
  clk, result, a, b
)/* synthesis syn_black_box syn_noprune=1 */;
  input clk;
  output [63 : 0] result;
  input [63 : 0] a;
  input [63 : 0] b;
  // synthesis translate_off
  wire sig00000001;
  wire sig00000002;
  wire sig00000003;
  wire sig00000004;
  wire sig00000005;
  wire sig00000006;
  wire sig00000007;
  wire sig00000008;
  wire sig00000009;
  wire sig0000000a;
  wire sig0000000b;
  wire sig0000000c;
  wire sig0000000d;
  wire sig0000000e;
  wire sig0000000f;
  wire sig00000010;
  wire sig00000011;
  wire sig00000012;
  wire sig00000013;
  wire sig00000014;
  wire sig00000015;
  wire sig00000016;
  wire sig00000017;
  wire sig00000018;
  wire sig00000019;
  wire sig0000001a;
  wire sig0000001b;
  wire sig0000001c;
  wire sig0000001d;
  wire sig0000001e;
  wire sig0000001f;
  wire sig00000020;
  wire sig00000021;
  wire sig00000022;
  wire sig00000023;
  wire sig00000024;
  wire sig00000025;
  wire sig00000026;
  wire sig00000027;
  wire sig00000028;
  wire sig00000029;
  wire sig0000002a;
  wire sig0000002b;
  wire sig0000002c;
  wire sig0000002d;
  wire sig0000002e;
  wire sig0000002f;
  wire sig00000030;
  wire sig00000031;
  wire sig00000032;
  wire sig00000033;
  wire sig00000034;
  wire sig00000035;
  wire sig00000036;
  wire sig00000037;
  wire sig00000038;
  wire sig00000039;
  wire sig0000003a;
  wire sig0000003b;
  wire sig0000003c;
  wire sig0000003d;
  wire sig0000003e;
  wire sig0000003f;
  wire sig00000040;
  wire sig00000041;
  wire sig00000042;
  wire sig00000043;
  wire sig00000044;
  wire sig00000045;
  wire sig00000046;
  wire sig00000047;
  wire sig00000048;
  wire sig00000049;
  wire sig0000004a;
  wire sig0000004b;
  wire sig0000004c;
  wire sig0000004d;
  wire sig0000004e;
  wire sig0000004f;
  wire sig00000050;
  wire sig00000051;
  wire sig00000052;
  wire sig00000053;
  wire sig00000054;
  wire sig00000055;
  wire sig00000056;
  wire sig00000057;
  wire sig00000058;
  wire sig00000059;
  wire sig0000005a;
  wire sig0000005b;
  wire sig0000005c;
  wire sig0000005d;
  wire sig0000005e;
  wire sig0000005f;
  wire sig00000060;
  wire sig00000061;
  wire sig00000062;
  wire sig00000063;
  wire sig00000064;
  wire sig00000065;
  wire sig00000066;
  wire sig00000067;
  wire sig00000068;
  wire sig00000069;
  wire sig0000006a;
  wire sig0000006b;
  wire sig0000006c;
  wire sig0000006d;
  wire sig0000006e;
  wire sig0000006f;
  wire sig00000070;
  wire sig00000071;
  wire sig00000072;
  wire sig00000073;
  wire sig00000074;
  wire sig00000075;
  wire sig00000076;
  wire sig00000077;
  wire sig00000078;
  wire sig00000079;
  wire sig0000007a;
  wire sig0000007b;
  wire sig0000007c;
  wire sig0000007d;
  wire sig0000007e;
  wire sig0000007f;
  wire sig00000080;
  wire sig00000081;
  wire sig00000082;
  wire sig00000083;
  wire sig00000084;
  wire sig00000085;
  wire sig00000086;
  wire sig00000087;
  wire sig00000088;
  wire sig00000089;
  wire sig0000008a;
  wire sig0000008b;
  wire sig0000008c;
  wire sig0000008d;
  wire sig0000008e;
  wire sig0000008f;
  wire sig00000090;
  wire sig00000091;
  wire sig00000092;
  wire sig00000093;
  wire sig00000094;
  wire sig00000095;
  wire sig00000096;
  wire sig00000097;
  wire sig00000098;
  wire sig00000099;
  wire sig0000009a;
  wire sig0000009b;
  wire sig0000009c;
  wire sig0000009d;
  wire sig0000009e;
  wire sig0000009f;
  wire sig000000a0;
  wire sig000000a1;
  wire sig000000a2;
  wire sig000000a3;
  wire sig000000a4;
  wire sig000000a5;
  wire sig000000a6;
  wire sig000000a7;
  wire sig000000a8;
  wire sig000000a9;
  wire sig000000aa;
  wire sig000000ab;
  wire sig000000ac;
  wire sig000000ad;
  wire sig000000ae;
  wire sig000000af;
  wire sig000000b0;
  wire sig000000b1;
  wire sig000000b2;
  wire sig000000b3;
  wire sig000000b4;
  wire sig000000b5;
  wire sig000000b6;
  wire sig000000b7;
  wire sig000000b8;
  wire sig000000b9;
  wire sig000000ba;
  wire sig000000bb;
  wire sig000000bc;
  wire sig000000bd;
  wire sig000000be;
  wire sig000000bf;
  wire sig000000c0;
  wire sig000000c1;
  wire sig000000c2;
  wire sig000000c3;
  wire sig000000c4;
  wire sig000000c5;
  wire sig000000c6;
  wire sig000000c7;
  wire sig000000c8;
  wire sig000000c9;
  wire sig000000ca;
  wire sig000000cb;
  wire sig000000cc;
  wire sig000000cd;
  wire sig000000ce;
  wire sig000000cf;
  wire sig000000d0;
  wire sig000000d1;
  wire sig000000d2;
  wire sig000000d3;
  wire sig000000d4;
  wire sig000000d5;
  wire sig000000d6;
  wire sig000000d7;
  wire sig000000d8;
  wire sig000000d9;
  wire sig000000da;
  wire sig000000db;
  wire sig000000dc;
  wire sig000000dd;
  wire sig000000de;
  wire sig000000df;
  wire sig000000e0;
  wire sig000000e1;
  wire sig000000e2;
  wire sig000000e3;
  wire sig000000e4;
  wire sig000000e5;
  wire sig000000e6;
  wire sig000000e7;
  wire sig000000e8;
  wire sig000000e9;
  wire sig000000ea;
  wire sig000000eb;
  wire sig000000ec;
  wire sig000000ed;
  wire sig000000ee;
  wire sig000000ef;
  wire sig000000f0;
  wire sig000000f1;
  wire sig000000f2;
  wire sig000000f3;
  wire sig000000f4;
  wire sig000000f5;
  wire sig000000f6;
  wire sig000000f7;
  wire sig000000f8;
  wire sig000000f9;
  wire sig000000fa;
  wire sig000000fb;
  wire sig000000fc;
  wire sig000000fd;
  wire sig000000fe;
  wire sig000000ff;
  wire sig00000100;
  wire sig00000101;
  wire sig00000102;
  wire sig00000103;
  wire sig00000104;
  wire sig00000105;
  wire sig00000106;
  wire sig00000107;
  wire sig00000108;
  wire sig00000109;
  wire sig0000010a;
  wire sig0000010b;
  wire sig0000010c;
  wire sig0000010d;
  wire sig0000010e;
  wire sig0000010f;
  wire sig00000110;
  wire sig00000111;
  wire sig00000112;
  wire sig00000113;
  wire sig00000114;
  wire sig00000115;
  wire sig00000116;
  wire sig00000117;
  wire sig00000118;
  wire sig00000119;
  wire sig0000011a;
  wire sig0000011b;
  wire sig0000011c;
  wire sig0000011d;
  wire sig0000011e;
  wire sig0000011f;
  wire sig00000120;
  wire sig00000121;
  wire sig00000122;
  wire sig00000123;
  wire sig00000124;
  wire sig00000125;
  wire sig00000126;
  wire sig00000127;
  wire sig00000128;
  wire sig00000129;
  wire sig0000012a;
  wire sig0000012b;
  wire sig0000012c;
  wire sig0000012d;
  wire sig0000012e;
  wire sig0000012f;
  wire sig00000130;
  wire sig00000131;
  wire sig00000132;
  wire sig00000133;
  wire sig00000134;
  wire sig00000135;
  wire sig00000136;
  wire sig00000137;
  wire sig00000138;
  wire sig00000139;
  wire sig0000013a;
  wire sig0000013b;
  wire sig0000013c;
  wire sig0000013d;
  wire sig0000013e;
  wire sig0000013f;
  wire sig00000140;
  wire sig00000141;
  wire sig00000142;
  wire sig00000143;
  wire sig00000144;
  wire sig00000145;
  wire sig00000146;
  wire sig00000147;
  wire sig00000148;
  wire sig00000149;
  wire sig0000014a;
  wire sig0000014b;
  wire sig0000014c;
  wire sig0000014d;
  wire sig0000014e;
  wire sig0000014f;
  wire sig00000150;
  wire sig00000151;
  wire sig00000152;
  wire sig00000153;
  wire sig00000154;
  wire sig00000155;
  wire sig00000156;
  wire sig00000157;
  wire sig00000158;
  wire sig00000159;
  wire sig0000015a;
  wire sig0000015b;
  wire sig0000015c;
  wire sig0000015d;
  wire sig0000015e;
  wire sig0000015f;
  wire sig00000160;
  wire sig00000161;
  wire sig00000162;
  wire sig00000163;
  wire sig00000164;
  wire sig00000165;
  wire sig00000166;
  wire sig00000167;
  wire sig00000168;
  wire sig00000169;
  wire sig0000016a;
  wire sig0000016b;
  wire sig0000016c;
  wire sig0000016d;
  wire sig0000016e;
  wire sig0000016f;
  wire sig00000170;
  wire sig00000171;
  wire sig00000172;
  wire sig00000173;
  wire sig00000174;
  wire sig00000175;
  wire sig00000176;
  wire sig00000177;
  wire sig00000178;
  wire sig00000179;
  wire sig0000017a;
  wire sig0000017b;
  wire sig0000017c;
  wire sig0000017d;
  wire sig0000017e;
  wire sig0000017f;
  wire sig00000180;
  wire sig00000181;
  wire sig00000182;
  wire sig00000183;
  wire sig00000184;
  wire sig00000185;
  wire sig00000186;
  wire sig00000187;
  wire sig00000188;
  wire sig00000189;
  wire sig0000018a;
  wire sig0000018b;
  wire sig0000018c;
  wire sig0000018d;
  wire sig0000018e;
  wire sig0000018f;
  wire sig00000190;
  wire sig00000191;
  wire sig00000192;
  wire sig00000193;
  wire sig00000194;
  wire sig00000195;
  wire sig00000196;
  wire sig00000197;
  wire sig00000198;
  wire sig00000199;
  wire sig0000019a;
  wire sig0000019b;
  wire sig0000019c;
  wire sig0000019d;
  wire sig0000019e;
  wire sig0000019f;
  wire sig000001a0;
  wire sig000001a1;
  wire sig000001a2;
  wire sig000001a3;
  wire sig000001a4;
  wire sig000001a5;
  wire sig000001a6;
  wire sig000001a7;
  wire sig000001a8;
  wire sig000001a9;
  wire sig000001aa;
  wire sig000001ab;
  wire sig000001ac;
  wire sig000001ad;
  wire sig000001ae;
  wire sig000001af;
  wire sig000001b0;
  wire sig000001b1;
  wire sig000001b2;
  wire sig000001b3;
  wire sig000001b4;
  wire sig000001b5;
  wire sig000001b6;
  wire sig000001b7;
  wire sig000001b8;
  wire sig000001b9;
  wire sig000001ba;
  wire sig000001bb;
  wire sig000001bc;
  wire sig000001bd;
  wire sig000001be;
  wire sig000001bf;
  wire sig000001c0;
  wire sig000001c1;
  wire sig000001c2;
  wire sig000001c3;
  wire sig000001c4;
  wire sig000001c5;
  wire sig000001c6;
  wire sig000001c7;
  wire sig000001c8;
  wire sig000001c9;
  wire sig000001ca;
  wire sig000001cb;
  wire sig000001cc;
  wire sig000001cd;
  wire sig000001ce;
  wire sig000001cf;
  wire sig000001d0;
  wire sig000001d1;
  wire sig000001d2;
  wire sig000001d3;
  wire sig000001d4;
  wire sig000001d5;
  wire sig000001d6;
  wire sig000001d7;
  wire sig000001d8;
  wire sig000001d9;
  wire sig000001da;
  wire sig000001db;
  wire sig000001dc;
  wire sig000001dd;
  wire sig000001de;
  wire sig000001df;
  wire sig000001e0;
  wire sig000001e1;
  wire sig000001e2;
  wire sig000001e3;
  wire sig000001e4;
  wire sig000001e5;
  wire sig000001e6;
  wire sig000001e7;
  wire sig000001e8;
  wire sig000001e9;
  wire sig000001ea;
  wire sig000001eb;
  wire sig000001ec;
  wire sig000001ed;
  wire sig000001ee;
  wire sig000001ef;
  wire sig000001f0;
  wire sig000001f1;
  wire sig000001f2;
  wire sig000001f3;
  wire sig000001f4;
  wire sig000001f5;
  wire sig000001f6;
  wire sig000001f7;
  wire sig000001f8;
  wire sig000001f9;
  wire sig000001fa;
  wire sig000001fb;
  wire sig000001fc;
  wire sig000001fd;
  wire sig000001fe;
  wire sig000001ff;
  wire sig00000200;
  wire sig00000201;
  wire sig00000202;
  wire sig00000203;
  wire sig00000204;
  wire sig00000205;
  wire sig00000206;
  wire sig00000207;
  wire sig00000208;
  wire sig00000209;
  wire sig0000020a;
  wire sig0000020b;
  wire sig0000020c;
  wire sig0000020d;
  wire sig0000020e;
  wire sig0000020f;
  wire sig00000210;
  wire sig00000211;
  wire sig00000212;
  wire sig00000213;
  wire sig00000214;
  wire sig00000215;
  wire sig00000216;
  wire sig00000217;
  wire sig00000218;
  wire sig00000219;
  wire sig0000021a;
  wire sig0000021b;
  wire sig0000021c;
  wire sig0000021d;
  wire sig0000021e;
  wire sig0000021f;
  wire sig00000220;
  wire sig00000221;
  wire sig00000222;
  wire sig00000223;
  wire sig00000224;
  wire sig00000225;
  wire sig00000226;
  wire sig00000227;
  wire sig00000228;
  wire sig00000229;
  wire sig0000022a;
  wire sig0000022b;
  wire sig0000022c;
  wire sig0000022d;
  wire sig0000022e;
  wire sig0000022f;
  wire sig00000230;
  wire sig00000231;
  wire sig00000232;
  wire sig00000233;
  wire sig00000234;
  wire sig00000235;
  wire sig00000236;
  wire sig00000237;
  wire sig00000238;
  wire sig00000239;
  wire sig0000023a;
  wire sig0000023b;
  wire sig0000023c;
  wire sig0000023d;
  wire sig0000023e;
  wire sig0000023f;
  wire sig00000240;
  wire sig00000241;
  wire sig00000242;
  wire sig00000243;
  wire sig00000244;
  wire sig00000245;
  wire sig00000246;
  wire sig00000247;
  wire sig00000248;
  wire sig00000249;
  wire sig0000024a;
  wire sig0000024b;
  wire sig0000024c;
  wire sig0000024d;
  wire sig0000024e;
  wire sig0000024f;
  wire sig00000250;
  wire sig00000251;
  wire sig00000252;
  wire sig00000253;
  wire sig00000254;
  wire sig00000255;
  wire sig00000256;
  wire sig00000257;
  wire sig00000258;
  wire sig00000259;
  wire sig0000025a;
  wire sig0000025b;
  wire sig0000025c;
  wire sig0000025d;
  wire sig0000025e;
  wire sig0000025f;
  wire sig00000260;
  wire sig00000261;
  wire sig00000262;
  wire sig00000263;
  wire sig00000264;
  wire sig00000265;
  wire sig00000266;
  wire sig00000267;
  wire sig00000268;
  wire sig00000269;
  wire sig0000026a;
  wire sig0000026b;
  wire sig0000026c;
  wire sig0000026d;
  wire sig0000026e;
  wire sig0000026f;
  wire sig00000270;
  wire sig00000271;
  wire sig00000272;
  wire sig00000273;
  wire sig00000274;
  wire sig00000275;
  wire sig00000276;
  wire sig00000277;
  wire sig00000278;
  wire sig00000279;
  wire sig0000027a;
  wire sig0000027b;
  wire sig0000027c;
  wire sig0000027d;
  wire sig0000027e;
  wire sig0000027f;
  wire sig00000280;
  wire sig00000281;
  wire sig00000282;
  wire sig00000283;
  wire sig00000284;
  wire sig00000285;
  wire sig00000286;
  wire sig00000287;
  wire sig00000288;
  wire sig00000289;
  wire sig0000028a;
  wire sig0000028b;
  wire sig0000028c;
  wire sig0000028d;
  wire sig0000028e;
  wire sig0000028f;
  wire sig00000290;
  wire sig00000291;
  wire sig00000292;
  wire sig00000293;
  wire sig00000294;
  wire sig00000295;
  wire sig00000296;
  wire sig00000297;
  wire sig00000298;
  wire sig00000299;
  wire sig0000029a;
  wire sig0000029b;
  wire sig0000029c;
  wire sig0000029d;
  wire sig0000029e;
  wire sig0000029f;
  wire sig000002a0;
  wire sig000002a1;
  wire sig000002a2;
  wire sig000002a3;
  wire sig000002a4;
  wire sig000002a5;
  wire sig000002a6;
  wire sig000002a7;
  wire sig000002a8;
  wire sig000002a9;
  wire sig000002aa;
  wire sig000002ab;
  wire sig000002ac;
  wire sig000002ad;
  wire sig000002ae;
  wire sig000002af;
  wire sig000002b0;
  wire sig000002b1;
  wire sig000002b2;
  wire sig000002b3;
  wire sig000002b4;
  wire sig000002b5;
  wire sig000002b6;
  wire sig000002b7;
  wire sig000002b8;
  wire sig000002b9;
  wire sig000002ba;
  wire sig000002bb;
  wire sig000002bc;
  wire sig000002bd;
  wire sig000002be;
  wire sig000002bf;
  wire sig000002c0;
  wire sig000002c1;
  wire sig000002c2;
  wire sig000002c3;
  wire sig000002c4;
  wire sig000002c5;
  wire sig000002c6;
  wire sig000002c7;
  wire sig000002c8;
  wire sig000002c9;
  wire sig000002ca;
  wire sig000002cb;
  wire sig000002cc;
  wire sig000002cd;
  wire sig000002ce;
  wire sig000002cf;
  wire sig000002d0;
  wire sig000002d1;
  wire sig000002d2;
  wire sig000002d3;
  wire sig000002d4;
  wire sig000002d5;
  wire sig000002d6;
  wire sig000002d7;
  wire sig000002d8;
  wire sig000002d9;
  wire sig000002da;
  wire sig000002db;
  wire sig000002dc;
  wire sig000002dd;
  wire sig000002de;
  wire sig000002df;
  wire sig000002e0;
  wire sig000002e1;
  wire sig000002e2;
  wire sig000002e3;
  wire sig000002e4;
  wire sig000002e5;
  wire sig000002e6;
  wire sig000002e7;
  wire sig000002e8;
  wire sig000002e9;
  wire sig000002ea;
  wire sig000002eb;
  wire sig000002ec;
  wire sig000002ed;
  wire sig000002ee;
  wire sig000002ef;
  wire sig000002f0;
  wire sig000002f1;
  wire sig000002f2;
  wire sig000002f3;
  wire sig000002f4;
  wire sig000002f5;
  wire sig000002f6;
  wire sig000002f7;
  wire sig000002f8;
  wire sig000002f9;
  wire sig000002fa;
  wire sig000002fb;
  wire sig000002fc;
  wire sig000002fd;
  wire sig000002fe;
  wire sig000002ff;
  wire sig00000300;
  wire sig00000301;
  wire sig00000302;
  wire sig00000303;
  wire sig00000304;
  wire sig00000305;
  wire sig00000306;
  wire sig00000307;
  wire sig00000308;
  wire sig00000309;
  wire sig0000030a;
  wire sig0000030b;
  wire sig0000030c;
  wire sig0000030d;
  wire sig0000030e;
  wire sig0000030f;
  wire sig00000310;
  wire sig00000311;
  wire sig00000312;
  wire sig00000313;
  wire sig00000314;
  wire sig00000315;
  wire sig00000316;
  wire sig00000317;
  wire sig00000318;
  wire sig00000319;
  wire sig0000031a;
  wire sig0000031b;
  wire sig0000031c;
  wire sig0000031d;
  wire sig0000031e;
  wire sig0000031f;
  wire sig00000320;
  wire sig00000321;
  wire sig00000322;
  wire sig00000323;
  wire sig00000324;
  wire sig00000325;
  wire sig00000326;
  wire sig00000327;
  wire sig00000328;
  wire sig00000329;
  wire sig0000032a;
  wire sig0000032b;
  wire sig0000032c;
  wire sig0000032d;
  wire sig0000032e;
  wire sig0000032f;
  wire sig00000330;
  wire sig00000331;
  wire sig00000332;
  wire sig00000333;
  wire sig00000334;
  wire sig00000335;
  wire sig00000336;
  wire sig00000337;
  wire sig00000338;
  wire sig00000339;
  wire sig0000033a;
  wire sig0000033b;
  wire sig0000033c;
  wire sig0000033d;
  wire sig0000033e;
  wire sig0000033f;
  wire sig00000340;
  wire sig00000341;
  wire sig00000342;
  wire sig00000343;
  wire sig00000344;
  wire sig00000345;
  wire sig00000346;
  wire sig00000347;
  wire sig00000348;
  wire sig00000349;
  wire sig0000034a;
  wire sig0000034b;
  wire sig0000034c;
  wire sig0000034d;
  wire sig0000034e;
  wire sig0000034f;
  wire sig00000350;
  wire sig00000351;
  wire sig00000352;
  wire sig00000353;
  wire sig00000354;
  wire sig00000355;
  wire sig00000356;
  wire sig00000357;
  wire sig00000358;
  wire sig00000359;
  wire sig0000035a;
  wire sig0000035b;
  wire sig0000035c;
  wire sig0000035d;
  wire sig0000035e;
  wire sig0000035f;
  wire sig00000360;
  wire sig00000361;
  wire sig00000362;
  wire sig00000363;
  wire sig00000364;
  wire sig00000365;
  wire sig00000366;
  wire sig00000367;
  wire sig00000368;
  wire sig00000369;
  wire sig0000036a;
  wire sig0000036b;
  wire sig0000036c;
  wire sig0000036d;
  wire sig0000036e;
  wire sig0000036f;
  wire sig00000370;
  wire sig00000371;
  wire sig00000372;
  wire sig00000373;
  wire sig00000374;
  wire sig00000375;
  wire sig00000376;
  wire sig00000377;
  wire sig00000378;
  wire sig00000379;
  wire sig0000037a;
  wire sig0000037b;
  wire sig0000037c;
  wire sig0000037d;
  wire sig0000037e;
  wire sig0000037f;
  wire sig00000380;
  wire sig00000381;
  wire sig00000382;
  wire sig00000383;
  wire sig00000384;
  wire sig00000385;
  wire sig00000386;
  wire sig00000387;
  wire sig00000388;
  wire sig00000389;
  wire sig0000038a;
  wire sig0000038b;
  wire sig0000038c;
  wire sig0000038d;
  wire sig0000038e;
  wire sig0000038f;
  wire sig00000390;
  wire sig00000391;
  wire sig00000392;
  wire sig00000393;
  wire sig00000394;
  wire sig00000395;
  wire sig00000396;
  wire sig00000397;
  wire sig00000398;
  wire sig00000399;
  wire sig0000039a;
  wire sig0000039b;
  wire sig0000039c;
  wire sig0000039d;
  wire sig0000039e;
  wire sig0000039f;
  wire sig000003a0;
  wire sig000003a1;
  wire sig000003a2;
  wire sig000003a3;
  wire sig000003a4;
  wire sig000003a5;
  wire sig000003a6;
  wire sig000003a7;
  wire sig000003a8;
  wire sig000003a9;
  wire sig000003aa;
  wire sig000003ab;
  wire sig000003ac;
  wire sig000003ad;
  wire sig000003ae;
  wire sig000003af;
  wire sig000003b0;
  wire sig000003b1;
  wire sig000003b2;
  wire sig000003b3;
  wire sig000003b4;
  wire sig000003b5;
  wire sig000003b6;
  wire sig000003b7;
  wire sig000003b8;
  wire sig000003b9;
  wire sig000003ba;
  wire sig000003bb;
  wire sig000003bc;
  wire sig000003bd;
  wire sig000003be;
  wire sig000003bf;
  wire sig000003c0;
  wire sig000003c1;
  wire sig000003c2;
  wire sig000003c3;
  wire sig000003c4;
  wire sig000003c5;
  wire sig000003c6;
  wire sig000003c7;
  wire sig000003c8;
  wire sig000003c9;
  wire sig000003ca;
  wire sig000003cb;
  wire sig000003cc;
  wire sig000003cd;
  wire sig000003ce;
  wire sig000003cf;
  wire sig000003d0;
  wire sig000003d1;
  wire sig000003d2;
  wire sig000003d3;
  wire sig000003d4;
  wire sig000003d5;
  wire sig000003d6;
  wire sig000003d7;
  wire sig000003d8;
  wire sig000003d9;
  wire sig000003da;
  wire sig000003db;
  wire sig000003dc;
  wire sig000003dd;
  wire sig000003de;
  wire sig000003df;
  wire sig000003e0;
  wire sig000003e1;
  wire sig000003e2;
  wire sig000003e3;
  wire sig000003e4;
  wire sig000003e5;
  wire sig000003e6;
  wire sig000003e7;
  wire sig000003e8;
  wire sig000003e9;
  wire sig000003ea;
  wire sig000003eb;
  wire sig000003ec;
  wire sig000003ed;
  wire sig000003ee;
  wire sig000003ef;
  wire sig000003f0;
  wire sig000003f1;
  wire sig000003f2;
  wire sig000003f3;
  wire sig000003f4;
  wire sig000003f5;
  wire sig000003f6;
  wire sig000003f7;
  wire sig000003f8;
  wire sig000003f9;
  wire sig000003fa;
  wire sig000003fb;
  wire sig000003fc;
  wire sig000003fd;
  wire sig000003fe;
  wire sig000003ff;
  wire sig00000400;
  wire sig00000401;
  wire sig00000402;
  wire sig00000403;
  wire sig00000404;
  wire sig00000405;
  wire sig00000406;
  wire sig00000407;
  wire sig00000408;
  wire sig00000409;
  wire sig0000040a;
  wire sig0000040b;
  wire sig0000040c;
  wire sig0000040d;
  wire sig0000040e;
  wire sig0000040f;
  wire sig00000410;
  wire sig00000411;
  wire sig00000412;
  wire sig00000413;
  wire sig00000414;
  wire sig00000415;
  wire sig00000416;
  wire sig00000417;
  wire sig00000418;
  wire sig00000419;
  wire sig0000041a;
  wire sig0000041b;
  wire sig0000041c;
  wire sig0000041d;
  wire sig0000041e;
  wire sig0000041f;
  wire sig00000420;
  wire sig00000421;
  wire sig00000422;
  wire sig00000423;
  wire sig00000424;
  wire sig00000425;
  wire sig00000426;
  wire sig00000427;
  wire sig00000428;
  wire sig00000429;
  wire sig0000042a;
  wire sig0000042b;
  wire sig0000042c;
  wire sig0000042d;
  wire sig0000042e;
  wire sig0000042f;
  wire sig00000430;
  wire sig00000431;
  wire sig00000432;
  wire sig00000433;
  wire sig00000434;
  wire sig00000435;
  wire sig00000436;
  wire sig00000437;
  wire sig00000438;
  wire sig00000439;
  wire sig0000043a;
  wire sig0000043b;
  wire sig0000043c;
  wire sig0000043d;
  wire sig0000043e;
  wire sig0000043f;
  wire sig00000440;
  wire sig00000441;
  wire sig00000442;
  wire sig00000443;
  wire sig00000444;
  wire sig00000445;
  wire sig00000446;
  wire sig00000447;
  wire sig00000448;
  wire sig00000449;
  wire sig0000044a;
  wire sig0000044b;
  wire sig0000044c;
  wire sig0000044d;
  wire sig0000044e;
  wire sig0000044f;
  wire sig00000450;
  wire sig00000451;
  wire sig00000452;
  wire sig00000453;
  wire sig00000454;
  wire sig00000455;
  wire sig00000456;
  wire sig00000457;
  wire sig00000458;
  wire sig00000459;
  wire sig0000045a;
  wire sig0000045b;
  wire sig0000045c;
  wire sig0000045d;
  wire sig0000045e;
  wire sig0000045f;
  wire sig00000460;
  wire sig00000461;
  wire sig00000462;
  wire sig00000463;
  wire sig00000464;
  wire sig00000465;
  wire sig00000466;
  wire sig00000467;
  wire sig00000468;
  wire sig00000469;
  wire sig0000046a;
  wire sig0000046b;
  wire sig0000046c;
  wire sig0000046d;
  wire sig0000046e;
  wire sig0000046f;
  wire sig00000470;
  wire sig00000471;
  wire sig00000472;
  wire sig00000473;
  wire sig00000474;
  wire sig00000475;
  wire sig00000476;
  wire sig00000477;
  wire sig00000478;
  wire sig00000479;
  wire sig0000047a;
  wire sig0000047b;
  wire sig0000047c;
  wire sig0000047d;
  wire sig0000047e;
  wire sig0000047f;
  wire sig00000480;
  wire sig00000481;
  wire sig00000482;
  wire sig00000483;
  wire sig00000484;
  wire sig00000485;
  wire sig00000486;
  wire sig00000487;
  wire sig00000488;
  wire sig00000489;
  wire sig0000048a;
  wire sig0000048b;
  wire sig0000048c;
  wire sig0000048d;
  wire sig0000048e;
  wire sig0000048f;
  wire sig00000490;
  wire sig00000491;
  wire sig00000492;
  wire sig00000493;
  wire sig00000494;
  wire sig00000495;
  wire sig00000496;
  wire sig00000497;
  wire sig00000498;
  wire sig00000499;
  wire sig0000049a;
  wire sig0000049b;
  wire sig0000049c;
  wire sig0000049d;
  wire sig0000049e;
  wire sig0000049f;
  wire sig000004a0;
  wire sig000004a1;
  wire sig000004a2;
  wire sig000004a3;
  wire sig000004a4;
  wire sig000004a5;
  wire sig000004a6;
  wire sig000004a7;
  wire sig000004a8;
  wire sig000004a9;
  wire sig000004aa;
  wire sig000004ab;
  wire sig000004ac;
  wire sig000004ad;
  wire sig000004ae;
  wire sig000004af;
  wire sig000004b0;
  wire sig000004b1;
  wire sig000004b2;
  wire sig000004b3;
  wire sig000004b4;
  wire sig000004b5;
  wire sig000004b6;
  wire sig000004b7;
  wire sig000004b8;
  wire sig000004b9;
  wire sig000004ba;
  wire sig000004bb;
  wire sig000004bc;
  wire sig000004bd;
  wire sig000004be;
  wire sig000004bf;
  wire sig000004c0;
  wire sig000004c1;
  wire sig000004c2;
  wire sig000004c3;
  wire sig000004c4;
  wire sig000004c5;
  wire sig000004c6;
  wire sig000004c7;
  wire sig000004c8;
  wire sig000004c9;
  wire sig000004ca;
  wire sig000004cb;
  wire sig000004cc;
  wire sig000004cd;
  wire sig000004ce;
  wire sig000004cf;
  wire sig000004d0;
  wire sig000004d1;
  wire sig000004d2;
  wire sig000004d3;
  wire sig000004d4;
  wire sig000004d5;
  wire sig000004d6;
  wire sig000004d7;
  wire sig000004d8;
  wire sig000004d9;
  wire sig000004da;
  wire sig000004db;
  wire sig000004dc;
  wire sig000004dd;
  wire sig000004de;
  wire sig000004df;
  wire sig000004e0;
  wire sig000004e1;
  wire sig000004e2;
  wire sig000004e3;
  wire sig000004e4;
  wire sig000004e5;
  wire sig000004e6;
  wire sig000004e7;
  wire sig000004e8;
  wire sig000004e9;
  wire sig000004ea;
  wire sig000004eb;
  wire sig000004ec;
  wire sig000004ed;
  wire sig000004ee;
  wire sig000004ef;
  wire sig000004f0;
  wire sig000004f1;
  wire sig000004f2;
  wire sig000004f3;
  wire sig000004f4;
  wire sig000004f5;
  wire sig000004f6;
  wire sig000004f7;
  wire sig000004f8;
  wire sig000004f9;
  wire sig000004fa;
  wire sig000004fb;
  wire sig000004fc;
  wire sig000004fd;
  wire sig000004fe;
  wire sig000004ff;
  wire sig00000500;
  wire sig00000501;
  wire sig00000502;
  wire sig00000503;
  wire sig00000504;
  wire sig00000505;
  wire sig00000506;
  wire sig00000507;
  wire sig00000508;
  wire sig00000509;
  wire sig0000050a;
  wire sig0000050b;
  wire sig0000050c;
  wire sig0000050d;
  wire sig0000050e;
  wire sig0000050f;
  wire sig00000510;
  wire sig00000511;
  wire sig00000512;
  wire sig00000513;
  wire sig00000514;
  wire sig00000515;
  wire sig00000516;
  wire sig00000517;
  wire sig00000518;
  wire sig00000519;
  wire sig0000051a;
  wire sig0000051b;
  wire sig0000051c;
  wire sig0000051d;
  wire sig0000051e;
  wire sig0000051f;
  wire sig00000520;
  wire sig00000521;
  wire sig00000522;
  wire sig00000523;
  wire sig00000524;
  wire sig00000525;
  wire sig00000526;
  wire sig00000527;
  wire sig00000528;
  wire sig00000529;
  wire sig0000052a;
  wire sig0000052b;
  wire sig0000052c;
  wire sig0000052d;
  wire sig0000052e;
  wire sig0000052f;
  wire sig00000530;
  wire sig00000531;
  wire sig00000532;
  wire sig00000533;
  wire sig00000534;
  wire sig00000535;
  wire sig00000536;
  wire sig00000537;
  wire sig00000538;
  wire sig00000539;
  wire sig0000053a;
  wire sig0000053b;
  wire sig0000053c;
  wire sig0000053d;
  wire sig0000053e;
  wire sig0000053f;
  wire sig00000540;
  wire sig00000541;
  wire sig00000542;
  wire sig00000543;
  wire sig00000544;
  wire sig00000545;
  wire sig00000546;
  wire sig00000547;
  wire sig00000548;
  wire sig00000549;
  wire sig0000054a;
  wire sig0000054b;
  wire sig0000054c;
  wire sig0000054d;
  wire sig0000054e;
  wire sig0000054f;
  wire sig00000550;
  wire sig00000551;
  wire sig00000552;
  wire sig00000553;
  wire sig00000554;
  wire sig00000555;
  wire sig00000556;
  wire sig00000557;
  wire sig00000558;
  wire sig00000559;
  wire sig0000055a;
  wire sig0000055b;
  wire sig0000055c;
  wire sig0000055d;
  wire sig0000055e;
  wire sig0000055f;
  wire sig00000560;
  wire sig00000561;
  wire sig00000562;
  wire sig00000563;
  wire sig00000564;
  wire sig00000565;
  wire sig00000566;
  wire sig00000567;
  wire sig00000568;
  wire sig00000569;
  wire sig0000056a;
  wire sig0000056b;
  wire sig0000056c;
  wire sig0000056d;
  wire sig0000056e;
  wire sig0000056f;
  wire sig00000570;
  wire sig00000571;
  wire sig00000572;
  wire sig00000573;
  wire sig00000574;
  wire sig00000575;
  wire sig00000576;
  wire sig00000577;
  wire sig00000578;
  wire sig00000579;
  wire sig0000057a;
  wire sig0000057b;
  wire sig0000057c;
  wire sig0000057d;
  wire sig0000057e;
  wire sig0000057f;
  wire sig00000580;
  wire sig00000581;
  wire sig00000582;
  wire sig00000583;
  wire sig00000584;
  wire sig00000585;
  wire sig00000586;
  wire sig00000587;
  wire sig00000588;
  wire sig00000589;
  wire sig0000058a;
  wire sig0000058b;
  wire sig0000058c;
  wire sig0000058d;
  wire sig0000058e;
  wire sig0000058f;
  wire sig00000590;
  wire sig00000591;
  wire sig00000592;
  wire sig00000593;
  wire sig00000594;
  wire sig00000595;
  wire sig00000596;
  wire sig00000597;
  wire sig00000598;
  wire sig00000599;
  wire sig0000059a;
  wire sig0000059b;
  wire sig0000059c;
  wire sig0000059d;
  wire sig0000059e;
  wire sig0000059f;
  wire sig000005a0;
  wire sig000005a1;
  wire sig000005a2;
  wire sig000005a3;
  wire sig000005a4;
  wire sig000005a5;
  wire sig000005a6;
  wire sig000005a7;
  wire sig000005a8;
  wire sig000005a9;
  wire sig000005aa;
  wire sig000005ab;
  wire sig000005ac;
  wire sig000005ad;
  wire sig000005ae;
  wire sig000005af;
  wire sig000005b0;
  wire sig000005b1;
  wire sig000005b2;
  wire sig000005b3;
  wire sig000005b4;
  wire sig000005b5;
  wire sig000005b6;
  wire sig000005b7;
  wire sig000005b8;
  wire sig000005b9;
  wire sig000005ba;
  wire sig000005bb;
  wire sig000005bc;
  wire sig000005bd;
  wire sig000005be;
  wire sig000005bf;
  wire sig000005c0;
  wire sig000005c1;
  wire sig000005c2;
  wire sig000005c3;
  wire sig000005c4;
  wire sig000005c5;
  wire sig000005c6;
  wire sig000005c7;
  wire sig000005c8;
  wire sig000005c9;
  wire sig000005ca;
  wire sig000005cb;
  wire sig000005cc;
  wire sig000005cd;
  wire sig000005ce;
  wire sig000005cf;
  wire sig000005d0;
  wire sig000005d1;
  wire sig000005d2;
  wire sig000005d3;
  wire sig000005d4;
  wire sig000005d5;
  wire sig000005d6;
  wire sig000005d7;
  wire sig000005d8;
  wire sig000005d9;
  wire sig000005da;
  wire sig000005db;
  wire sig000005dc;
  wire sig000005dd;
  wire sig000005de;
  wire sig000005df;
  wire sig000005e0;
  wire sig000005e1;
  wire sig000005e2;
  wire sig000005e3;
  wire sig000005e4;
  wire sig000005e5;
  wire sig000005e6;
  wire sig000005e7;
  wire sig000005e8;
  wire sig000005e9;
  wire sig000005ea;
  wire sig000005eb;
  wire sig000005ec;
  wire sig000005ed;
  wire sig000005ee;
  wire sig000005ef;
  wire sig000005f0;
  wire sig000005f1;
  wire sig000005f2;
  wire sig000005f3;
  wire sig000005f4;
  wire sig000005f5;
  wire sig000005f6;
  wire sig000005f7;
  wire sig000005f8;
  wire sig000005f9;
  wire sig000005fa;
  wire sig000005fb;
  wire sig000005fc;
  wire sig000005fd;
  wire sig000005fe;
  wire sig000005ff;
  wire sig00000600;
  wire sig00000601;
  wire sig00000602;
  wire sig00000603;
  wire sig00000604;
  wire sig00000605;
  wire sig00000606;
  wire sig00000607;
  wire sig00000608;
  wire sig00000609;
  wire sig0000060a;
  wire sig0000060b;
  wire sig0000060c;
  wire sig0000060d;
  wire sig0000060e;
  wire sig0000060f;
  wire sig00000610;
  wire sig00000611;
  wire sig00000612;
  wire sig00000613;
  wire sig00000614;
  wire sig00000615;
  wire sig00000616;
  wire sig00000617;
  wire sig00000618;
  wire sig00000619;
  wire sig0000061a;
  wire sig0000061b;
  wire sig0000061c;
  wire sig0000061d;
  wire sig0000061e;
  wire sig0000061f;
  wire sig00000620;
  wire sig00000621;
  wire sig00000622;
  wire sig00000623;
  wire sig00000624;
  wire sig00000625;
  wire sig00000626;
  wire sig00000627;
  wire sig00000628;
  wire sig00000629;
  wire sig0000062a;
  wire sig0000062b;
  wire sig0000062c;
  wire sig0000062d;
  wire sig0000062e;
  wire sig0000062f;
  wire sig00000630;
  wire sig00000631;
  wire sig00000632;
  wire sig00000633;
  wire sig00000634;
  wire sig00000635;
  wire sig00000636;
  wire sig00000637;
  wire sig00000638;
  wire sig00000639;
  wire sig0000063a;
  wire sig0000063b;
  wire sig0000063c;
  wire sig0000063d;
  wire sig0000063e;
  wire sig0000063f;
  wire sig00000640;
  wire sig00000641;
  wire sig00000642;
  wire sig00000643;
  wire sig00000644;
  wire sig00000645;
  wire sig00000646;
  wire sig00000647;
  wire sig00000648;
  wire sig00000649;
  wire sig0000064a;
  wire sig0000064b;
  wire sig0000064c;
  wire sig0000064d;
  wire sig0000064e;
  wire sig0000064f;
  wire sig00000650;
  wire sig00000651;
  wire sig00000652;
  wire sig00000653;
  wire sig00000654;
  wire sig00000655;
  wire sig00000656;
  wire sig00000657;
  wire sig00000658;
  wire sig00000659;
  wire sig0000065a;
  wire sig0000065b;
  wire sig0000065c;
  wire sig0000065d;
  wire sig0000065e;
  wire sig0000065f;
  wire sig00000660;
  wire sig00000661;
  wire sig00000662;
  wire sig00000663;
  wire sig00000664;
  wire sig00000665;
  wire sig00000666;
  wire sig00000667;
  wire sig00000668;
  wire sig00000669;
  wire sig0000066a;
  wire sig0000066b;
  wire sig0000066c;
  wire sig0000066d;
  wire sig0000066e;
  wire sig0000066f;
  wire sig00000670;
  wire sig00000671;
  wire sig00000672;
  wire sig00000673;
  wire sig00000674;
  wire sig00000675;
  wire sig00000676;
  wire sig00000677;
  wire sig00000678;
  wire sig00000679;
  wire sig0000067a;
  wire sig0000067b;
  wire sig0000067c;
  wire sig0000067d;
  wire sig0000067e;
  wire sig0000067f;
  wire sig00000680;
  wire sig00000681;
  wire sig00000682;
  wire sig00000683;
  wire sig00000684;
  wire sig00000685;
  wire sig00000686;
  wire sig00000687;
  wire sig00000688;
  wire sig00000689;
  wire sig0000068a;
  wire sig0000068b;
  wire sig0000068c;
  wire sig0000068d;
  wire sig0000068e;
  wire sig0000068f;
  wire sig00000690;
  wire sig00000691;
  wire sig00000692;
  wire sig00000693;
  wire sig00000694;
  wire sig00000695;
  wire sig00000696;
  wire sig00000697;
  wire sig00000698;
  wire sig00000699;
  wire sig0000069a;
  wire sig0000069b;
  wire sig0000069c;
  wire sig0000069d;
  wire sig0000069e;
  wire sig0000069f;
  wire sig000006a0;
  wire sig000006a1;
  wire sig000006a2;
  wire sig000006a3;
  wire sig000006a4;
  wire sig000006a5;
  wire sig000006a6;
  wire sig000006a7;
  wire sig000006a8;
  wire sig000006a9;
  wire sig000006aa;
  wire sig000006ab;
  wire sig000006ac;
  wire sig000006ad;
  wire sig000006ae;
  wire sig000006af;
  wire sig000006b0;
  wire sig000006b1;
  wire sig000006b2;
  wire sig000006b3;
  wire sig000006b4;
  wire sig000006b5;
  wire sig000006b6;
  wire sig000006b7;
  wire sig000006b8;
  wire sig000006b9;
  wire sig000006ba;
  wire sig000006bb;
  wire sig000006bc;
  wire sig000006bd;
  wire sig000006be;
  wire sig000006bf;
  wire sig000006c0;
  wire sig000006c1;
  wire sig000006c2;
  wire sig000006c3;
  wire sig000006c4;
  wire sig000006c5;
  wire sig000006c6;
  wire sig000006c7;
  wire sig000006c8;
  wire sig000006c9;
  wire sig000006ca;
  wire sig000006cb;
  wire sig000006cc;
  wire sig000006cd;
  wire sig000006ce;
  wire sig000006cf;
  wire sig000006d0;
  wire sig000006d1;
  wire sig000006d2;
  wire sig000006d3;
  wire sig000006d4;
  wire sig000006d5;
  wire sig000006d6;
  wire sig000006d7;
  wire sig000006d8;
  wire sig000006d9;
  wire sig000006da;
  wire sig000006db;
  wire sig000006dc;
  wire sig000006dd;
  wire sig000006de;
  wire sig000006df;
  wire sig000006e0;
  wire sig000006e1;
  wire sig000006e2;
  wire sig000006e3;
  wire sig000006e4;
  wire sig000006e5;
  wire sig000006e6;
  wire sig000006e7;
  wire sig000006e8;
  wire sig000006e9;
  wire sig000006ea;
  wire sig000006eb;
  wire sig000006ec;
  wire sig000006ed;
  wire sig000006ee;
  wire sig000006ef;
  wire sig000006f0;
  wire sig000006f1;
  wire sig000006f2;
  wire sig000006f3;
  wire sig000006f4;
  wire sig000006f5;
  wire sig000006f6;
  wire sig000006f7;
  wire sig000006f8;
  wire sig000006f9;
  wire sig000006fa;
  wire sig000006fb;
  wire sig000006fc;
  wire sig000006fd;
  wire sig000006fe;
  wire sig000006ff;
  wire sig00000700;
  wire sig00000701;
  wire sig00000702;
  wire sig00000703;
  wire sig00000704;
  wire sig00000705;
  wire sig00000706;
  wire sig00000707;
  wire sig00000708;
  wire sig00000709;
  wire sig0000070a;
  wire sig0000070b;
  wire sig0000070c;
  wire sig0000070d;
  wire sig0000070e;
  wire sig0000070f;
  wire sig00000710;
  wire sig00000711;
  wire sig00000712;
  wire sig00000713;
  wire sig00000714;
  wire sig00000715;
  wire sig00000716;
  wire sig00000717;
  wire sig00000718;
  wire sig00000719;
  wire sig0000071a;
  wire sig0000071b;
  wire sig0000071c;
  wire sig0000071d;
  wire sig0000071e;
  wire sig0000071f;
  wire sig00000720;
  wire sig00000721;
  wire sig00000722;
  wire sig00000723;
  wire sig00000724;
  wire sig00000725;
  wire sig00000726;
  wire sig00000727;
  wire sig00000728;
  wire sig00000729;
  wire sig0000072a;
  wire sig0000072b;
  wire sig0000072c;
  wire sig0000072d;
  wire sig0000072e;
  wire sig0000072f;
  wire sig00000730;
  wire sig00000731;
  wire sig00000732;
  wire sig00000733;
  wire sig00000734;
  wire sig00000735;
  wire sig00000736;
  wire sig00000737;
  wire sig00000738;
  wire sig00000739;
  wire sig0000073a;
  wire sig0000073b;
  wire sig0000073c;
  wire sig0000073d;
  wire sig0000073e;
  wire sig0000073f;
  wire sig00000740;
  wire sig00000741;
  wire sig00000742;
  wire sig00000743;
  wire sig00000744;
  wire sig00000745;
  wire sig00000746;
  wire sig00000747;
  wire sig00000748;
  wire sig00000749;
  wire sig0000074a;
  wire sig0000074b;
  wire sig0000074c;
  wire sig0000074d;
  wire sig0000074e;
  wire sig0000074f;
  wire sig00000750;
  wire sig00000751;
  wire sig00000752;
  wire sig00000753;
  wire sig00000754;
  wire sig00000755;
  wire sig00000756;
  wire sig00000757;
  wire sig00000758;
  wire sig00000759;
  wire sig0000075a;
  wire sig0000075b;
  wire sig0000075c;
  wire sig0000075d;
  wire sig0000075e;
  wire sig0000075f;
  wire sig00000760;
  wire sig00000761;
  wire sig00000762;
  wire sig00000763;
  wire sig00000764;
  wire sig00000765;
  wire sig00000766;
  wire sig00000767;
  wire sig00000768;
  wire sig00000769;
  wire sig0000076a;
  wire sig0000076b;
  wire sig0000076c;
  wire sig0000076d;
  wire sig0000076e;
  wire sig0000076f;
  wire sig00000770;
  wire sig00000771;
  wire sig00000772;
  wire sig00000773;
  wire sig00000774;
  wire sig00000775;
  wire sig00000776;
  wire sig00000777;
  wire sig00000778;
  wire sig00000779;
  wire sig0000077a;
  wire sig0000077b;
  wire sig0000077c;
  wire sig0000077d;
  wire sig0000077e;
  wire sig0000077f;
  wire sig00000780;
  wire sig00000781;
  wire sig00000782;
  wire sig00000783;
  wire sig00000784;
  wire sig00000785;
  wire sig00000786;
  wire sig00000787;
  wire sig00000788;
  wire sig00000789;
  wire sig0000078a;
  wire sig0000078b;
  wire sig0000078c;
  wire sig0000078d;
  wire sig0000078e;
  wire sig0000078f;
  wire sig00000790;
  wire sig00000791;
  wire sig00000792;
  wire sig00000793;
  wire sig00000794;
  wire sig00000795;
  wire sig00000796;
  wire sig00000797;
  wire sig00000798;
  wire sig00000799;
  wire sig0000079a;
  wire sig0000079b;
  wire sig0000079c;
  wire sig0000079d;
  wire sig0000079e;
  wire sig0000079f;
  wire sig000007a0;
  wire sig000007a1;
  wire sig000007a2;
  wire sig000007a3;
  wire sig000007a4;
  wire sig000007a5;
  wire sig000007a6;
  wire sig000007a7;
  wire sig000007a8;
  wire sig000007a9;
  wire sig000007aa;
  wire sig000007ab;
  wire sig000007ac;
  wire sig000007ad;
  wire sig000007ae;
  wire sig000007af;
  wire sig000007b0;
  wire sig000007b1;
  wire sig000007b2;
  wire sig000007b3;
  wire sig000007b4;
  wire sig000007b5;
  wire sig000007b6;
  wire sig000007b7;
  wire sig000007b8;
  wire sig000007b9;
  wire sig000007ba;
  wire sig000007bb;
  wire sig000007bc;
  wire sig000007bd;
  wire sig000007be;
  wire sig000007bf;
  wire sig000007c0;
  wire sig000007c1;
  wire sig000007c2;
  wire sig000007c3;
  wire sig000007c4;
  wire sig000007c5;
  wire sig000007c6;
  wire sig000007c7;
  wire sig000007c8;
  wire sig000007c9;
  wire sig000007ca;
  wire sig000007cb;
  wire sig000007cc;
  wire sig000007cd;
  wire sig000007ce;
  wire sig000007cf;
  wire sig000007d0;
  wire sig000007d1;
  wire sig000007d2;
  wire sig000007d3;
  wire sig000007d4;
  wire sig000007d5;
  wire sig000007d6;
  wire sig000007d7;
  wire sig000007d8;
  wire sig000007d9;
  wire sig000007da;
  wire sig000007db;
  wire sig000007dc;
  wire sig000007dd;
  wire sig000007de;
  wire sig000007df;
  wire sig000007e0;
  wire sig000007e1;
  wire sig000007e2;
  wire sig000007e3;
  wire sig000007e4;
  wire sig000007e5;
  wire sig000007e6;
  wire sig000007e7;
  wire sig000007e8;
  wire sig000007e9;
  wire sig000007ea;
  wire sig000007eb;
  wire sig000007ec;
  wire sig000007ed;
  wire sig000007ee;
  wire sig000007ef;
  wire sig000007f0;
  wire sig000007f1;
  wire sig000007f2;
  wire sig000007f3;
  wire sig000007f4;
  wire sig000007f5;
  wire sig000007f6;
  wire sig000007f7;
  wire sig000007f8;
  wire sig000007f9;
  wire sig000007fa;
  wire sig000007fb;
  wire sig000007fc;
  wire sig000007fd;
  wire sig000007fe;
  wire sig000007ff;
  wire sig00000800;
  wire sig00000801;
  wire sig00000802;
  wire sig00000803;
  wire sig00000804;
  wire sig00000805;
  wire sig00000806;
  wire sig00000807;
  wire sig00000808;
  wire sig00000809;
  wire sig0000080a;
  wire sig0000080b;
  wire sig0000080c;
  wire sig0000080d;
  wire sig0000080e;
  wire sig0000080f;
  wire sig00000810;
  wire sig00000811;
  wire sig00000812;
  wire sig00000813;
  wire sig00000814;
  wire sig00000815;
  wire sig00000816;
  wire sig00000817;
  wire sig00000818;
  wire sig00000819;
  wire sig0000081a;
  wire sig0000081b;
  wire sig0000081c;
  wire sig0000081d;
  wire sig0000081e;
  wire sig0000081f;
  wire sig00000820;
  wire sig00000821;
  wire sig00000822;
  wire sig00000823;
  wire sig00000824;
  wire sig00000825;
  wire sig00000826;
  wire sig00000827;
  wire sig00000828;
  wire sig00000829;
  wire sig0000082a;
  wire sig0000082b;
  wire sig0000082c;
  wire sig0000082d;
  wire sig0000082e;
  wire sig0000082f;
  wire sig00000830;
  wire sig00000831;
  wire sig00000832;
  wire sig00000833;
  wire sig00000834;
  wire sig00000835;
  wire sig00000836;
  wire sig00000837;
  wire sig00000838;
  wire sig00000839;
  wire sig0000083a;
  wire sig0000083b;
  wire sig0000083c;
  wire sig0000083d;
  wire sig0000083e;
  wire sig0000083f;
  wire sig00000840;
  wire sig00000841;
  wire sig00000842;
  wire sig00000843;
  wire sig00000844;
  wire sig00000845;
  wire sig00000846;
  wire sig00000847;
  wire sig00000848;
  wire sig00000849;
  wire sig0000084a;
  wire sig0000084b;
  wire sig0000084c;
  wire sig0000084d;
  wire sig0000084e;
  wire sig0000084f;
  wire sig00000850;
  wire sig00000851;
  wire sig00000852;
  wire sig00000853;
  wire sig00000854;
  wire sig00000855;
  wire sig00000856;
  wire sig00000857;
  wire sig00000858;
  wire sig00000859;
  wire sig0000085a;
  wire sig0000085b;
  wire sig0000085c;
  wire sig0000085d;
  wire sig0000085e;
  wire sig0000085f;
  wire sig00000860;
  wire sig00000861;
  wire sig00000862;
  wire sig00000863;
  wire sig00000864;
  wire sig00000865;
  wire sig00000866;
  wire sig00000867;
  wire sig00000868;
  wire sig00000869;
  wire sig0000086a;
  wire sig0000086b;
  wire sig0000086c;
  wire sig0000086d;
  wire sig0000086e;
  wire sig0000086f;
  wire sig00000870;
  wire sig00000871;
  wire sig00000872;
  wire sig00000873;
  wire sig00000874;
  wire sig00000875;
  wire sig00000876;
  wire sig00000877;
  wire sig00000878;
  wire sig00000879;
  wire sig0000087a;
  wire sig0000087b;
  wire sig0000087c;
  wire sig0000087d;
  wire sig0000087e;
  wire sig0000087f;
  wire sig00000880;
  wire sig00000881;
  wire sig00000882;
  wire sig00000883;
  wire sig00000884;
  wire sig00000885;
  wire sig00000886;
  wire sig00000887;
  wire sig00000888;
  wire sig00000889;
  wire sig0000088a;
  wire sig0000088b;
  wire sig0000088c;
  wire sig0000088d;
  wire sig0000088e;
  wire sig0000088f;
  wire sig00000890;
  wire sig00000891;
  wire sig00000892;
  wire sig00000893;
  wire sig00000894;
  wire sig00000895;
  wire sig00000896;
  wire sig00000897;
  wire sig00000898;
  wire sig00000899;
  wire sig0000089a;
  wire sig0000089b;
  wire sig0000089c;
  wire sig0000089d;
  wire sig0000089e;
  wire sig0000089f;
  wire sig000008a0;
  wire sig000008a1;
  wire sig000008a2;
  wire sig000008a3;
  wire sig000008a4;
  wire sig000008a5;
  wire sig000008a6;
  wire sig000008a7;
  wire sig000008a8;
  wire sig000008a9;
  wire sig000008aa;
  wire sig000008ab;
  wire sig000008ac;
  wire sig000008ad;
  wire sig000008ae;
  wire sig000008af;
  wire sig000008b0;
  wire sig000008b1;
  wire sig000008b2;
  wire sig000008b3;
  wire sig000008b4;
  wire sig000008b5;
  wire sig000008b6;
  wire sig000008b7;
  wire sig000008b8;
  wire \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op ;
  wire sig000008b9;
  wire sig000008ba;
  wire sig000008bb;
  wire sig000008bc;
  wire NLW_blk000002f9_O_UNCONNECTED;
  wire NLW_blk000002fa_O_UNCONNECTED;
  wire NLW_blk000002fc_O_UNCONNECTED;
  wire NLW_blk000002fe_O_UNCONNECTED;
  wire NLW_blk00000300_O_UNCONNECTED;
  wire NLW_blk00000302_O_UNCONNECTED;
  wire NLW_blk00000304_O_UNCONNECTED;
  wire NLW_blk00000306_O_UNCONNECTED;
  wire NLW_blk00000308_O_UNCONNECTED;
  wire NLW_blk0000030a_O_UNCONNECTED;
  wire NLW_blk0000030c_O_UNCONNECTED;
  wire NLW_blk000003d9_O_UNCONNECTED;
  wire NLW_blk00000875_Q15_UNCONNECTED;
  wire NLW_blk00000877_Q15_UNCONNECTED;
  wire NLW_blk00000879_Q15_UNCONNECTED;
  wire NLW_blk0000087b_Q15_UNCONNECTED;
  wire NLW_blk0000087d_Q15_UNCONNECTED;
  wire NLW_blk0000087f_Q15_UNCONNECTED;
  wire NLW_blk00000881_Q15_UNCONNECTED;
  wire NLW_blk00000883_Q15_UNCONNECTED;
  wire NLW_blk00000885_Q15_UNCONNECTED;
  wire NLW_blk00000887_Q15_UNCONNECTED;
  wire NLW_blk00000889_Q15_UNCONNECTED;
  wire NLW_blk0000088b_Q15_UNCONNECTED;
  wire NLW_blk0000088d_Q15_UNCONNECTED;
  wire NLW_blk0000088f_Q15_UNCONNECTED;
  wire NLW_blk00000891_Q15_UNCONNECTED;
  wire NLW_blk00000893_Q15_UNCONNECTED;
  wire NLW_blk00000895_Q15_UNCONNECTED;
  wire NLW_blk00000897_Q15_UNCONNECTED;
  wire NLW_blk00000899_Q15_UNCONNECTED;
  wire NLW_blk0000089b_Q15_UNCONNECTED;
  wire NLW_blk0000089d_Q15_UNCONNECTED;
  wire NLW_blk0000089f_Q15_UNCONNECTED;
  wire NLW_blk000008a1_Q15_UNCONNECTED;
  wire NLW_blk000008a3_Q15_UNCONNECTED;
  wire NLW_blk000008a5_Q15_UNCONNECTED;
  wire NLW_blk000008a7_Q15_UNCONNECTED;
  wire NLW_blk000008a9_Q15_UNCONNECTED;
  wire NLW_blk000008ab_Q15_UNCONNECTED;
  wire NLW_blk000008ad_Q15_UNCONNECTED;
  wire NLW_blk000008af_Q15_UNCONNECTED;
  wire NLW_blk000008b1_Q15_UNCONNECTED;
  wire NLW_blk000008b3_Q15_UNCONNECTED;
  wire NLW_blk000008b5_Q15_UNCONNECTED;
  wire NLW_blk000008b7_Q15_UNCONNECTED;
  wire NLW_blk000008b9_Q15_UNCONNECTED;
  wire NLW_blk000008bb_Q15_UNCONNECTED;
  wire NLW_blk000008bd_Q15_UNCONNECTED;
  wire NLW_blk000008bf_Q15_UNCONNECTED;
  wire NLW_blk000008c1_Q15_UNCONNECTED;
  wire NLW_blk000008c3_Q15_UNCONNECTED;
  wire NLW_blk000008c5_Q15_UNCONNECTED;
  wire NLW_blk000008c7_Q15_UNCONNECTED;
  wire NLW_blk000008c9_Q15_UNCONNECTED;
  wire NLW_blk000008cb_Q15_UNCONNECTED;
  wire NLW_blk000008cd_Q15_UNCONNECTED;
  wire NLW_blk000008cf_Q15_UNCONNECTED;
  wire NLW_blk000008d1_Q15_UNCONNECTED;
  wire NLW_blk000008d3_Q15_UNCONNECTED;
  wire NLW_blk000008d5_Q15_UNCONNECTED;
  wire NLW_blk000008d7_Q15_UNCONNECTED;
  wire NLW_blk000008d9_Q15_UNCONNECTED;
  wire NLW_blk000008db_Q15_UNCONNECTED;
  wire NLW_blk000008dd_Q15_UNCONNECTED;
  wire NLW_blk000008df_Q15_UNCONNECTED;
  wire NLW_blk000008e1_Q15_UNCONNECTED;
  wire NLW_blk000008e3_Q15_UNCONNECTED;
  wire NLW_blk000008e5_Q15_UNCONNECTED;
  wire NLW_blk000008e7_Q15_UNCONNECTED;
  wire NLW_blk000008e9_Q15_UNCONNECTED;
  wire NLW_blk000008eb_Q15_UNCONNECTED;
  wire NLW_blk000008ed_Q15_UNCONNECTED;
  wire NLW_blk000008ef_Q15_UNCONNECTED;
  wire NLW_blk000008f1_Q15_UNCONNECTED;
  wire NLW_blk000008f3_Q15_UNCONNECTED;
  wire NLW_blk000008f5_Q15_UNCONNECTED;
  wire NLW_blk000008f7_Q15_UNCONNECTED;
  wire NLW_blk000008f9_Q15_UNCONNECTED;
  wire NLW_blk000008fb_Q15_UNCONNECTED;
  wire NLW_blk000008fd_Q15_UNCONNECTED;
  wire NLW_blk000008ff_Q15_UNCONNECTED;
  wire NLW_blk00000901_Q15_UNCONNECTED;
  wire NLW_blk00000903_Q15_UNCONNECTED;
  wire NLW_blk00000905_Q15_UNCONNECTED;
  wire NLW_blk00000907_Q15_UNCONNECTED;
  wire [10 : 0] \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op ;
  wire [51 : 0] \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op ;
  assign
    result[63] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op ,
    result[62] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [10],
    result[61] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [9],
    result[60] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [8],
    result[59] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [7],
    result[58] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [6],
    result[57] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [5],
    result[56] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [4],
    result[55] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [3],
    result[54] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [2],
    result[53] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [1],
    result[52] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [0],
    result[51] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [51],
    result[50] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [50],
    result[49] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [49],
    result[48] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [48],
    result[47] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [47],
    result[46] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [46],
    result[45] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [45],
    result[44] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [44],
    result[43] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [43],
    result[42] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [42],
    result[41] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [41],
    result[40] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [40],
    result[39] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [39],
    result[38] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [38],
    result[37] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [37],
    result[36] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [36],
    result[35] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [35],
    result[34] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [34],
    result[33] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [33],
    result[32] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [32],
    result[31] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [31],
    result[30] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [30],
    result[29] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [29],
    result[28] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [28],
    result[27] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [27],
    result[26] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [26],
    result[25] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [25],
    result[24] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [24],
    result[23] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [23],
    result[22] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [22],
    result[21] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [21],
    result[20] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [20],
    result[19] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [19],
    result[18] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [18],
    result[17] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [17],
    result[16] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [16],
    result[15] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [15],
    result[14] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [14],
    result[13] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [13],
    result[12] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [12],
    result[11] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [11],
    result[10] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [10],
    result[9] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [9],
    result[8] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [8],
    result[7] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [7],
    result[6] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [6],
    result[5] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [5],
    result[4] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [4],
    result[3] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [3],
    result[2] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [2],
    result[1] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [1],
    result[0] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [0];
  GND   blk00000001 (
    .G(sig00000001)
  );
  VCC   blk00000002 (
    .P(sig00000002)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000003 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000003df),
    .Q(sig0000035e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000004 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000003dd),
    .Q(sig0000035a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000005 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000130),
    .Q(sig0000035b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000006 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000035c),
    .Q(sig0000035d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000007 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000008bc),
    .Q(sig0000035c)
  );
  MUXCY   blk00000008 (
    .CI(sig00000001),
    .DI(sig00000458),
    .S(sig00000316),
    .O(sig00000315)
  );
  XORCY   blk00000009 (
    .CI(sig00000001),
    .LI(sig00000316),
    .O(sig00000369)
  );
  MUXCY   blk0000000a (
    .CI(sig00000315),
    .DI(sig00000001),
    .S(sig00000360),
    .O(sig00000317)
  );
  XORCY   blk0000000b (
    .CI(sig00000315),
    .LI(sig00000360),
    .O(sig0000036b)
  );
  MUXCY   blk0000000c (
    .CI(sig00000317),
    .DI(sig00000001),
    .S(sig00000361),
    .O(sig00000318)
  );
  XORCY   blk0000000d (
    .CI(sig00000317),
    .LI(sig00000361),
    .O(sig0000036c)
  );
  MUXCY   blk0000000e (
    .CI(sig00000318),
    .DI(sig00000001),
    .S(sig00000362),
    .O(sig00000319)
  );
  XORCY   blk0000000f (
    .CI(sig00000318),
    .LI(sig00000362),
    .O(sig0000036d)
  );
  MUXCY   blk00000010 (
    .CI(sig00000319),
    .DI(sig00000001),
    .S(sig00000363),
    .O(sig0000031a)
  );
  XORCY   blk00000011 (
    .CI(sig00000319),
    .LI(sig00000363),
    .O(sig0000036e)
  );
  MUXCY   blk00000012 (
    .CI(sig0000031a),
    .DI(sig00000001),
    .S(sig00000364),
    .O(sig0000031b)
  );
  XORCY   blk00000013 (
    .CI(sig0000031a),
    .LI(sig00000364),
    .O(sig0000036f)
  );
  MUXCY   blk00000014 (
    .CI(sig0000031b),
    .DI(sig00000001),
    .S(sig00000365),
    .O(sig0000031c)
  );
  XORCY   blk00000015 (
    .CI(sig0000031b),
    .LI(sig00000365),
    .O(sig00000370)
  );
  MUXCY   blk00000016 (
    .CI(sig0000031c),
    .DI(sig00000001),
    .S(sig00000366),
    .O(sig0000031d)
  );
  XORCY   blk00000017 (
    .CI(sig0000031c),
    .LI(sig00000366),
    .O(sig00000371)
  );
  MUXCY   blk00000018 (
    .CI(sig0000031d),
    .DI(sig00000001),
    .S(sig00000367),
    .O(sig0000031e)
  );
  XORCY   blk00000019 (
    .CI(sig0000031d),
    .LI(sig00000367),
    .O(sig00000372)
  );
  MUXCY   blk0000001a (
    .CI(sig0000031e),
    .DI(sig00000001),
    .S(sig00000368),
    .O(sig0000031f)
  );
  XORCY   blk0000001b (
    .CI(sig0000031e),
    .LI(sig00000368),
    .O(sig00000373)
  );
  XORCY   blk0000001c (
    .CI(sig0000031f),
    .LI(sig0000035f),
    .O(sig0000036a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000001d (
    .C(clk),
    .D(sig000003d6),
    .Q(sig0000034f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000001e (
    .C(clk),
    .D(sig000003d5),
    .Q(sig0000034e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000001f (
    .C(clk),
    .D(sig000003d3),
    .Q(sig0000034c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000020 (
    .C(clk),
    .D(sig000003d2),
    .Q(sig0000034b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000021 (
    .C(clk),
    .D(sig000003d1),
    .Q(sig0000034a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000022 (
    .C(clk),
    .D(sig000003d0),
    .Q(sig00000349)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000023 (
    .C(clk),
    .D(sig000003cf),
    .Q(sig00000348)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000024 (
    .C(clk),
    .D(sig000003ce),
    .Q(sig00000347)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000025 (
    .C(clk),
    .D(sig000003cd),
    .Q(sig00000346)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000026 (
    .C(clk),
    .D(sig000003cc),
    .Q(sig00000345)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000027 (
    .C(clk),
    .D(sig000003cb),
    .Q(sig00000344)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000028 (
    .C(clk),
    .D(sig000003ca),
    .Q(sig00000343)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000029 (
    .C(clk),
    .D(sig000003c8),
    .Q(sig00000341)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000002a (
    .C(clk),
    .D(sig000003c7),
    .Q(sig00000340)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000002b (
    .C(clk),
    .D(sig000003c6),
    .Q(sig0000033f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000002c (
    .C(clk),
    .D(sig000003c5),
    .Q(sig0000033e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000002d (
    .C(clk),
    .D(sig000003c4),
    .Q(sig0000033d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000002e (
    .C(clk),
    .D(sig000003c3),
    .Q(sig0000033c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000002f (
    .C(clk),
    .D(sig000003c2),
    .Q(sig0000033b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000030 (
    .C(clk),
    .D(sig000003c1),
    .Q(sig0000033a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000031 (
    .C(clk),
    .D(sig000003c0),
    .Q(sig00000339)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000032 (
    .C(clk),
    .D(sig000003bf),
    .Q(sig00000338)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000033 (
    .C(clk),
    .D(sig000003bd),
    .Q(sig00000336)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000034 (
    .C(clk),
    .D(sig000003bc),
    .Q(sig00000335)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000035 (
    .C(clk),
    .D(sig000003bb),
    .Q(sig00000334)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000036 (
    .C(clk),
    .D(sig000003ba),
    .Q(sig00000333)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000037 (
    .C(clk),
    .D(sig000003b9),
    .Q(sig00000332)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000038 (
    .C(clk),
    .D(sig000003b8),
    .Q(sig00000331)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000039 (
    .C(clk),
    .D(sig000003b7),
    .Q(sig00000330)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000003a (
    .C(clk),
    .D(sig000003b6),
    .Q(sig0000032f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000003b (
    .C(clk),
    .D(sig000003b5),
    .Q(sig0000032e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000003c (
    .C(clk),
    .D(sig000003b4),
    .Q(sig0000032d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000003d (
    .C(clk),
    .D(sig000003b2),
    .Q(sig0000032b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000003e (
    .C(clk),
    .D(sig000003b1),
    .Q(sig0000032a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000003f (
    .C(clk),
    .D(sig000003b0),
    .Q(sig00000329)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000040 (
    .C(clk),
    .D(sig000003af),
    .Q(sig00000328)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000041 (
    .C(clk),
    .D(sig000003ae),
    .Q(sig00000327)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000042 (
    .C(clk),
    .D(sig000003ad),
    .Q(sig00000326)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000043 (
    .C(clk),
    .D(sig000003ac),
    .Q(sig00000325)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000044 (
    .C(clk),
    .D(sig000003ab),
    .Q(sig00000324)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000045 (
    .C(clk),
    .D(sig000003aa),
    .Q(sig00000323)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000046 (
    .C(clk),
    .D(sig000003a9),
    .Q(sig00000322)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000047 (
    .C(clk),
    .D(sig000003dc),
    .Q(sig00000355)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000048 (
    .C(clk),
    .D(sig000003db),
    .Q(sig00000354)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000049 (
    .C(clk),
    .D(sig000003da),
    .Q(sig00000353)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000004a (
    .C(clk),
    .D(sig000003d9),
    .Q(sig00000352)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000004b (
    .C(clk),
    .D(sig000003d8),
    .Q(sig0000034d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000004c (
    .C(clk),
    .D(sig000003d4),
    .Q(sig00000342)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000004d (
    .C(clk),
    .D(sig000003c9),
    .Q(sig00000337)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000004e (
    .C(clk),
    .D(sig000003be),
    .Q(sig0000032c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000004f (
    .C(clk),
    .D(sig000003b3),
    .Q(sig00000321)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000050 (
    .C(clk),
    .D(sig000003a8),
    .Q(sig00000320)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000051 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000036a),
    .Q(sig0000001e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000052 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000373),
    .Q(sig00000026)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000053 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000372),
    .Q(sig00000025)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000054 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000371),
    .Q(sig00000024)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000055 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000370),
    .Q(sig00000023)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000056 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000036f),
    .Q(sig00000022)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000057 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000036e),
    .Q(sig00000021)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000058 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000036d),
    .Q(sig00000020)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000059 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000036c),
    .Q(sig0000001f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005a (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000036b),
    .Q(sig0000001d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005b (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000369),
    .Q(sig0000001c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005c (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ce),
    .Q(sig00000027)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005d (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d9),
    .Q(sig00000028)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005e (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e4),
    .Q(sig00000033)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005f (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ef),
    .Q(sig0000003e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000060 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000fa),
    .Q(sig00000049)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000061 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000100),
    .Q(sig00000054)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000062 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000101),
    .Q(sig0000005a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000063 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000102),
    .Q(sig0000005b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000064 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000103),
    .Q(sig0000005c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000065 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000104),
    .Q(sig0000005d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000066 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000cf),
    .Q(sig00000029)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000067 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d0),
    .Q(sig0000002a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000068 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d1),
    .Q(sig0000002b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000069 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d2),
    .Q(sig0000002c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006a (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d3),
    .Q(sig0000002d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006b (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d4),
    .Q(sig0000002e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006c (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d5),
    .Q(sig0000002f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006d (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d6),
    .Q(sig00000030)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006e (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d7),
    .Q(sig00000031)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006f (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000d8),
    .Q(sig00000032)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000070 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000da),
    .Q(sig00000034)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000071 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000db),
    .Q(sig00000035)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000072 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000dc),
    .Q(sig00000036)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000073 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000dd),
    .Q(sig00000037)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000074 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000de),
    .Q(sig00000038)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000075 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000df),
    .Q(sig00000039)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000076 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e0),
    .Q(sig0000003a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000077 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e1),
    .Q(sig0000003b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000078 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e2),
    .Q(sig0000003c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000079 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e3),
    .Q(sig0000003d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007a (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e5),
    .Q(sig0000003f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007b (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e6),
    .Q(sig00000040)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007c (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e7),
    .Q(sig00000041)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007d (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e8),
    .Q(sig00000042)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007e (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000e9),
    .Q(sig00000043)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007f (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ea),
    .Q(sig00000044)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000080 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000eb),
    .Q(sig00000045)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000081 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ec),
    .Q(sig00000046)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000082 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ed),
    .Q(sig00000047)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000083 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ee),
    .Q(sig00000048)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000084 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f0),
    .Q(sig0000004a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000085 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f1),
    .Q(sig0000004b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000086 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f2),
    .Q(sig0000004c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000087 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f3),
    .Q(sig0000004d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000088 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f4),
    .Q(sig0000004e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000089 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f5),
    .Q(sig0000004f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008a (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f6),
    .Q(sig00000050)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008b (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f7),
    .Q(sig00000051)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008c (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f8),
    .Q(sig00000052)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008d (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000f9),
    .Q(sig00000053)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008e (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000fb),
    .Q(sig00000055)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008f (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000fc),
    .Q(sig00000056)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000090 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000fd),
    .Q(sig00000057)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000091 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000fe),
    .Q(sig00000058)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000092 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ff),
    .Q(sig00000059)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000093 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000097),
    .Q(sig0000005e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000094 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a2),
    .Q(sig0000005f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000095 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ad),
    .Q(sig0000006a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000096 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b8),
    .Q(sig00000075)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000097 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c3),
    .Q(sig00000080)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000098 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c9),
    .Q(sig0000008b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000099 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ca),
    .Q(sig00000091)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009a (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000cb),
    .Q(sig00000092)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009b (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000cc),
    .Q(sig00000093)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009c (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000cd),
    .Q(sig00000094)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009d (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000098),
    .Q(sig00000060)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009e (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000099),
    .Q(sig00000061)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009f (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000009a),
    .Q(sig00000062)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000009b),
    .Q(sig00000063)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000009c),
    .Q(sig00000064)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000009d),
    .Q(sig00000065)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000009e),
    .Q(sig00000066)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000009f),
    .Q(sig00000067)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a0),
    .Q(sig00000068)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a1),
    .Q(sig00000069)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a3),
    .Q(sig0000006b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a4),
    .Q(sig0000006c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a5),
    .Q(sig0000006d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000aa (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a6),
    .Q(sig0000006e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ab (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a7),
    .Q(sig0000006f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ac (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a8),
    .Q(sig00000070)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ad (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000a9),
    .Q(sig00000071)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ae (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000aa),
    .Q(sig00000072)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000af (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ab),
    .Q(sig00000073)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ac),
    .Q(sig00000074)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ae),
    .Q(sig00000076)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000af),
    .Q(sig00000077)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b0),
    .Q(sig00000078)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b1),
    .Q(sig00000079)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b2),
    .Q(sig0000007a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b3),
    .Q(sig0000007b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b4),
    .Q(sig0000007c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b5),
    .Q(sig0000007d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b6),
    .Q(sig0000007e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ba (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b7),
    .Q(sig0000007f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bb (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000b9),
    .Q(sig00000081)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bc (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000ba),
    .Q(sig00000082)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bd (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000bb),
    .Q(sig00000083)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000be (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000bc),
    .Q(sig00000084)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bf (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000bd),
    .Q(sig00000085)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000be),
    .Q(sig00000086)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000bf),
    .Q(sig00000087)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c0),
    .Q(sig00000088)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c1),
    .Q(sig00000089)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c2),
    .Q(sig0000008a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c4),
    .Q(sig0000008c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c5),
    .Q(sig0000008d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c6),
    .Q(sig0000008e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c7),
    .Q(sig0000008f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000000c8),
    .Q(sig00000090)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ca (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000001f),
    .Q(sig00000095)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cb (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000020),
    .Q(sig00000096)
  );
  MUXCY   blk000000cc (
    .CI(sig00000108),
    .DI(sig00000001),
    .S(sig00000117),
    .O(sig00000109)
  );
  MUXCY   blk000000cd (
    .CI(sig00000107),
    .DI(sig00000001),
    .S(sig00000116),
    .O(sig00000108)
  );
  MUXCY   blk000000ce (
    .CI(sig00000106),
    .DI(sig00000001),
    .S(sig00000115),
    .O(sig00000107)
  );
  MUXCY   blk000000cf (
    .CI(sig00000105),
    .DI(sig00000001),
    .S(sig00000114),
    .O(sig00000106)
  );
  MUXCY   blk000000d0 (
    .CI(sig00000112),
    .DI(sig00000001),
    .S(sig00000120),
    .O(sig00000105)
  );
  MUXCY   blk000000d1 (
    .CI(sig00000111),
    .DI(sig00000001),
    .S(sig0000011f),
    .O(sig00000112)
  );
  MUXCY   blk000000d2 (
    .CI(sig00000110),
    .DI(sig00000001),
    .S(sig0000011e),
    .O(sig00000111)
  );
  MUXCY   blk000000d3 (
    .CI(sig0000010f),
    .DI(sig00000001),
    .S(sig0000011d),
    .O(sig00000110)
  );
  MUXCY   blk000000d4 (
    .CI(sig0000010e),
    .DI(sig00000001),
    .S(sig0000011c),
    .O(sig0000010f)
  );
  MUXCY   blk000000d5 (
    .CI(sig0000010d),
    .DI(sig00000001),
    .S(sig0000011b),
    .O(sig0000010e)
  );
  MUXCY   blk000000d6 (
    .CI(sig0000010c),
    .DI(sig00000001),
    .S(sig0000011a),
    .O(sig0000010d)
  );
  MUXCY   blk000000d7 (
    .CI(sig0000010b),
    .DI(sig00000001),
    .S(sig00000119),
    .O(sig0000010c)
  );
  MUXCY   blk000000d8 (
    .CI(sig0000010a),
    .DI(sig00000001),
    .S(sig00000118),
    .O(sig0000010b)
  );
  MUXCY   blk000000d9 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000113),
    .O(sig0000010a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000da (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000109),
    .Q(sig00000139)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000db (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000108),
    .Q(sig00000138)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000dc (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000107),
    .Q(sig00000137)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000dd (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000106),
    .Q(sig00000136)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000de (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000105),
    .Q(sig00000135)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000df (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000112),
    .Q(sig00000142)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000111),
    .Q(sig00000141)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000110),
    .Q(sig00000140)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000010f),
    .Q(sig0000013f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000010e),
    .Q(sig0000013e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000010d),
    .Q(sig0000013d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000010c),
    .Q(sig0000013c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000010b),
    .Q(sig0000013b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000010a),
    .Q(sig0000013a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000143),
    .Q(sig00000121)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000148),
    .Q(sig00000122)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ea (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000149),
    .Q(sig00000128)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000eb (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000014a),
    .Q(sig00000129)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ec (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000014b),
    .Q(sig0000012a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ed (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000014c),
    .Q(sig0000012b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ee (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000014d),
    .Q(sig0000012c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ef (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000014e),
    .Q(sig0000012d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000014f),
    .Q(sig0000012e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000150),
    .Q(sig0000012f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000144),
    .Q(sig00000123)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000145),
    .Q(sig00000124)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000146),
    .Q(sig00000125)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000147),
    .Q(sig00000126)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000002),
    .Q(sig00000127)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000155),
    .Q(sig00000130)
  );
  MUXF8   blk000000f8 (
    .I0(sig00000133),
    .I1(sig00000134),
    .S(sig00000132),
    .O(sig00000155)
  );
  MUXF7   blk000000f9 (
    .I0(sig00000153),
    .I1(sig00000154),
    .S(sig00000131),
    .O(sig00000134)
  );
  MUXF7   blk000000fa (
    .I0(sig00000151),
    .I1(sig00000152),
    .S(sig00000131),
    .O(sig00000133)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fb (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000021),
    .Q(sig00000131)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fc (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000022),
    .Q(sig00000132)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fd (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000263),
    .Q(sig000002c0)
  );
  MUXCY   blk000000fe (
    .CI(sig000002bf),
    .DI(sig00000001),
    .S(sig000002c1),
    .O(sig00000252)
  );
  XORCY   blk000000ff (
    .CI(sig000002bf),
    .LI(sig000002c1),
    .O(sig00000264)
  );
  MUXCY   blk00000100 (
    .CI(sig00000252),
    .DI(sig00000001),
    .S(sig000002c2),
    .O(sig0000025b)
  );
  XORCY   blk00000101 (
    .CI(sig00000252),
    .LI(sig000002c2),
    .O(sig0000026f)
  );
  MUXCY   blk00000102 (
    .CI(sig0000025b),
    .DI(sig000001c4),
    .S(sig000002f2),
    .O(sig0000025c)
  );
  XORCY   blk00000103 (
    .CI(sig0000025b),
    .LI(sig000002f2),
    .O(sig00000277)
  );
  MUXCY   blk00000104 (
    .CI(sig0000025c),
    .DI(sig000001c5),
    .S(sig000002f3),
    .O(sig0000025d)
  );
  XORCY   blk00000105 (
    .CI(sig0000025c),
    .LI(sig000002f3),
    .O(sig00000278)
  );
  MUXCY   blk00000106 (
    .CI(sig0000025d),
    .DI(sig000001d0),
    .S(sig000002f4),
    .O(sig0000025e)
  );
  XORCY   blk00000107 (
    .CI(sig0000025d),
    .LI(sig000002f4),
    .O(sig00000279)
  );
  MUXCY   blk00000108 (
    .CI(sig0000025e),
    .DI(sig000001d6),
    .S(sig000002f5),
    .O(sig0000025f)
  );
  XORCY   blk00000109 (
    .CI(sig0000025e),
    .LI(sig000002f5),
    .O(sig0000027a)
  );
  MUXCY   blk0000010a (
    .CI(sig0000025f),
    .DI(sig000001d7),
    .S(sig000002f6),
    .O(sig00000260)
  );
  XORCY   blk0000010b (
    .CI(sig0000025f),
    .LI(sig000002f6),
    .O(sig0000027b)
  );
  MUXCY   blk0000010c (
    .CI(sig00000260),
    .DI(sig000001d8),
    .S(sig000002f7),
    .O(sig00000261)
  );
  XORCY   blk0000010d (
    .CI(sig00000260),
    .LI(sig000002f7),
    .O(sig0000027c)
  );
  MUXCY   blk0000010e (
    .CI(sig00000261),
    .DI(sig000001d9),
    .S(sig000002f8),
    .O(sig00000262)
  );
  XORCY   blk0000010f (
    .CI(sig00000261),
    .LI(sig000002f8),
    .O(sig0000027d)
  );
  MUXCY   blk00000110 (
    .CI(sig00000262),
    .DI(sig000001da),
    .S(sig000002e0),
    .O(sig00000248)
  );
  XORCY   blk00000111 (
    .CI(sig00000262),
    .LI(sig000002e0),
    .O(sig0000027e)
  );
  MUXCY   blk00000112 (
    .CI(sig00000248),
    .DI(sig000001db),
    .S(sig000002e1),
    .O(sig00000249)
  );
  XORCY   blk00000113 (
    .CI(sig00000248),
    .LI(sig000002e1),
    .O(sig00000265)
  );
  MUXCY   blk00000114 (
    .CI(sig00000249),
    .DI(sig000001dc),
    .S(sig000002e2),
    .O(sig0000024a)
  );
  XORCY   blk00000115 (
    .CI(sig00000249),
    .LI(sig000002e2),
    .O(sig00000266)
  );
  MUXCY   blk00000116 (
    .CI(sig0000024a),
    .DI(sig000001c6),
    .S(sig000002e3),
    .O(sig0000024b)
  );
  XORCY   blk00000117 (
    .CI(sig0000024a),
    .LI(sig000002e3),
    .O(sig00000267)
  );
  MUXCY   blk00000118 (
    .CI(sig0000024b),
    .DI(sig000001c7),
    .S(sig000002e4),
    .O(sig0000024c)
  );
  XORCY   blk00000119 (
    .CI(sig0000024b),
    .LI(sig000002e4),
    .O(sig00000268)
  );
  MUXCY   blk0000011a (
    .CI(sig0000024c),
    .DI(sig000001c8),
    .S(sig000002e5),
    .O(sig0000024d)
  );
  XORCY   blk0000011b (
    .CI(sig0000024c),
    .LI(sig000002e5),
    .O(sig00000269)
  );
  MUXCY   blk0000011c (
    .CI(sig0000024d),
    .DI(sig000001c9),
    .S(sig000002e6),
    .O(sig0000024e)
  );
  XORCY   blk0000011d (
    .CI(sig0000024d),
    .LI(sig000002e6),
    .O(sig0000026a)
  );
  MUXCY   blk0000011e (
    .CI(sig0000024e),
    .DI(sig000001ca),
    .S(sig000002e7),
    .O(sig0000024f)
  );
  XORCY   blk0000011f (
    .CI(sig0000024e),
    .LI(sig000002e7),
    .O(sig0000026b)
  );
  MUXCY   blk00000120 (
    .CI(sig0000024f),
    .DI(sig000001cb),
    .S(sig000002e8),
    .O(sig00000250)
  );
  XORCY   blk00000121 (
    .CI(sig0000024f),
    .LI(sig000002e8),
    .O(sig0000026c)
  );
  MUXCY   blk00000122 (
    .CI(sig00000250),
    .DI(sig000001cc),
    .S(sig000002e9),
    .O(sig00000251)
  );
  XORCY   blk00000123 (
    .CI(sig00000250),
    .LI(sig000002e9),
    .O(sig0000026d)
  );
  MUXCY   blk00000124 (
    .CI(sig00000251),
    .DI(sig000001cd),
    .S(sig000002ea),
    .O(sig00000253)
  );
  XORCY   blk00000125 (
    .CI(sig00000251),
    .LI(sig000002ea),
    .O(sig0000026e)
  );
  MUXCY   blk00000126 (
    .CI(sig00000253),
    .DI(sig000001ce),
    .S(sig000002eb),
    .O(sig00000254)
  );
  XORCY   blk00000127 (
    .CI(sig00000253),
    .LI(sig000002eb),
    .O(sig00000270)
  );
  MUXCY   blk00000128 (
    .CI(sig00000254),
    .DI(sig000001cf),
    .S(sig000002ec),
    .O(sig00000255)
  );
  XORCY   blk00000129 (
    .CI(sig00000254),
    .LI(sig000002ec),
    .O(sig00000271)
  );
  MUXCY   blk0000012a (
    .CI(sig00000255),
    .DI(sig000001d1),
    .S(sig000002ed),
    .O(sig00000256)
  );
  XORCY   blk0000012b (
    .CI(sig00000255),
    .LI(sig000002ed),
    .O(sig00000272)
  );
  MUXCY   blk0000012c (
    .CI(sig00000256),
    .DI(sig000001d2),
    .S(sig000002ee),
    .O(sig00000257)
  );
  XORCY   blk0000012d (
    .CI(sig00000256),
    .LI(sig000002ee),
    .O(sig00000273)
  );
  MUXCY   blk0000012e (
    .CI(sig00000257),
    .DI(sig000001d3),
    .S(sig000002ef),
    .O(sig00000258)
  );
  XORCY   blk0000012f (
    .CI(sig00000257),
    .LI(sig000002ef),
    .O(sig00000274)
  );
  MUXCY   blk00000130 (
    .CI(sig00000258),
    .DI(sig000001d4),
    .S(sig000002f0),
    .O(sig00000259)
  );
  XORCY   blk00000131 (
    .CI(sig00000258),
    .LI(sig000002f0),
    .O(sig00000275)
  );
  MUXCY   blk00000132 (
    .CI(sig00000259),
    .DI(sig000001d5),
    .S(sig000002f1),
    .O(sig0000025a)
  );
  XORCY   blk00000133 (
    .CI(sig00000259),
    .LI(sig000002f1),
    .O(sig00000276)
  );
  XORCY   blk00000134 (
    .CI(sig0000025a),
    .LI(sig00000001),
    .O(sig00000263)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000135 (
    .C(clk),
    .D(sig00000240),
    .Q(sig00000225)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000136 (
    .C(clk),
    .D(sig0000023f),
    .Q(sig00000224)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000137 (
    .C(clk),
    .D(sig0000023e),
    .Q(sig00000223)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000138 (
    .C(clk),
    .D(sig0000023d),
    .Q(sig00000222)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000139 (
    .C(clk),
    .D(sig0000023c),
    .Q(sig00000221)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000013a (
    .C(clk),
    .D(sig0000023b),
    .Q(sig00000220)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000013b (
    .C(clk),
    .D(sig0000023a),
    .Q(sig0000021f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000013c (
    .C(clk),
    .D(sig00000238),
    .Q(sig0000021d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000013d (
    .C(clk),
    .D(sig00000237),
    .Q(sig0000021c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000013e (
    .C(clk),
    .D(sig00000236),
    .Q(sig0000021b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000013f (
    .C(clk),
    .D(sig00000235),
    .Q(sig0000021a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000140 (
    .C(clk),
    .D(sig00000234),
    .Q(sig00000219)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000141 (
    .C(clk),
    .D(sig00000233),
    .Q(sig00000218)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000142 (
    .C(clk),
    .D(sig00000232),
    .Q(sig00000217)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000143 (
    .C(clk),
    .D(sig00000231),
    .Q(sig00000216)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000144 (
    .C(clk),
    .D(sig00000230),
    .Q(sig00000215)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000145 (
    .C(clk),
    .D(sig0000022f),
    .Q(sig00000214)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000146 (
    .C(clk),
    .D(sig00000247),
    .Q(sig0000022c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000147 (
    .C(clk),
    .D(sig00000246),
    .Q(sig0000022b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000148 (
    .C(clk),
    .D(sig00000245),
    .Q(sig0000022a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000149 (
    .C(clk),
    .D(sig00000244),
    .Q(sig00000229)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000014a (
    .C(clk),
    .D(sig00000243),
    .Q(sig00000228)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000014b (
    .C(clk),
    .D(sig00000242),
    .Q(sig00000227)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000014c (
    .C(clk),
    .D(sig00000241),
    .Q(sig00000226)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000014d (
    .C(clk),
    .D(sig00000239),
    .Q(sig0000021e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000014e (
    .C(clk),
    .D(sig0000022e),
    .Q(sig00000213)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000014f (
    .C(clk),
    .D(sig0000022d),
    .Q(sig00000212)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000150 (
    .C(clk),
    .D(sig00000276),
    .Q(sig00000240)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000151 (
    .C(clk),
    .D(sig00000275),
    .Q(sig0000023f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000152 (
    .C(clk),
    .D(sig00000274),
    .Q(sig0000023e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000153 (
    .C(clk),
    .D(sig00000273),
    .Q(sig0000023d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000154 (
    .C(clk),
    .D(sig00000272),
    .Q(sig0000023c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000155 (
    .C(clk),
    .D(sig00000271),
    .Q(sig0000023b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000156 (
    .C(clk),
    .D(sig00000270),
    .Q(sig0000023a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000157 (
    .C(clk),
    .D(sig0000026e),
    .Q(sig00000238)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000158 (
    .C(clk),
    .D(sig0000026d),
    .Q(sig00000237)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000159 (
    .C(clk),
    .D(sig0000026c),
    .Q(sig00000236)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000015a (
    .C(clk),
    .D(sig0000026b),
    .Q(sig00000235)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000015b (
    .C(clk),
    .D(sig0000026a),
    .Q(sig00000234)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000015c (
    .C(clk),
    .D(sig00000269),
    .Q(sig00000233)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000015d (
    .C(clk),
    .D(sig00000268),
    .Q(sig00000232)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000015e (
    .C(clk),
    .D(sig00000267),
    .Q(sig00000231)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000015f (
    .C(clk),
    .D(sig00000266),
    .Q(sig00000230)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000160 (
    .C(clk),
    .D(sig00000265),
    .Q(sig0000022f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000161 (
    .C(clk),
    .D(sig0000027e),
    .Q(sig00000247)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000162 (
    .C(clk),
    .D(sig0000027d),
    .Q(sig00000246)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000163 (
    .C(clk),
    .D(sig0000027c),
    .Q(sig00000245)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000164 (
    .C(clk),
    .D(sig0000027b),
    .Q(sig00000244)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000165 (
    .C(clk),
    .D(sig0000027a),
    .Q(sig00000243)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000166 (
    .C(clk),
    .D(sig00000279),
    .Q(sig00000242)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000167 (
    .C(clk),
    .D(sig00000278),
    .Q(sig00000241)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000168 (
    .C(clk),
    .D(sig00000277),
    .Q(sig00000239)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000169 (
    .C(clk),
    .D(sig0000026f),
    .Q(sig0000022e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000016a (
    .C(clk),
    .D(sig00000264),
    .Q(sig0000022d)
  );
  MUXCY   blk0000016b (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000281),
    .O(sig00000282)
  );
  MUXCY   blk0000016c (
    .CI(sig00000282),
    .DI(sig0000018f),
    .S(sig000002f9),
    .O(sig0000028d)
  );
  XORCY   blk0000016d (
    .CI(sig00000282),
    .LI(sig000002f9),
    .O(sig000002c3)
  );
  MUXCY   blk0000016e (
    .CI(sig0000028d),
    .DI(sig00000190),
    .S(sig00000304),
    .O(sig00000297)
  );
  XORCY   blk0000016f (
    .CI(sig0000028d),
    .LI(sig00000304),
    .O(sig000002ce)
  );
  MUXCY   blk00000170 (
    .CI(sig00000297),
    .DI(sig0000019b),
    .S(sig0000030d),
    .O(sig00000298)
  );
  XORCY   blk00000171 (
    .CI(sig00000297),
    .LI(sig0000030d),
    .O(sig000002d8)
  );
  MUXCY   blk00000172 (
    .CI(sig00000298),
    .DI(sig000001a4),
    .S(sig0000030e),
    .O(sig00000299)
  );
  XORCY   blk00000173 (
    .CI(sig00000298),
    .LI(sig0000030e),
    .O(sig000002d9)
  );
  MUXCY   blk00000174 (
    .CI(sig00000299),
    .DI(sig000001a5),
    .S(sig0000030f),
    .O(sig0000029a)
  );
  XORCY   blk00000175 (
    .CI(sig00000299),
    .LI(sig0000030f),
    .O(sig000002da)
  );
  MUXCY   blk00000176 (
    .CI(sig0000029a),
    .DI(sig000001a6),
    .S(sig00000310),
    .O(sig0000029b)
  );
  XORCY   blk00000177 (
    .CI(sig0000029a),
    .LI(sig00000310),
    .O(sig000002db)
  );
  MUXCY   blk00000178 (
    .CI(sig0000029b),
    .DI(sig000001a7),
    .S(sig00000311),
    .O(sig0000029c)
  );
  XORCY   blk00000179 (
    .CI(sig0000029b),
    .LI(sig00000311),
    .O(sig000002dc)
  );
  MUXCY   blk0000017a (
    .CI(sig0000029c),
    .DI(sig000001a8),
    .S(sig00000312),
    .O(sig0000029d)
  );
  XORCY   blk0000017b (
    .CI(sig0000029c),
    .LI(sig00000312),
    .O(sig000002dd)
  );
  MUXCY   blk0000017c (
    .CI(sig0000029d),
    .DI(sig000001a9),
    .S(sig00000313),
    .O(sig0000029e)
  );
  XORCY   blk0000017d (
    .CI(sig0000029d),
    .LI(sig00000313),
    .O(sig000002de)
  );
  MUXCY   blk0000017e (
    .CI(sig0000029e),
    .DI(sig000001aa),
    .S(sig00000314),
    .O(sig00000283)
  );
  XORCY   blk0000017f (
    .CI(sig0000029e),
    .LI(sig00000314),
    .O(sig000002df)
  );
  MUXCY   blk00000180 (
    .CI(sig00000283),
    .DI(sig00000191),
    .S(sig000002fa),
    .O(sig00000284)
  );
  XORCY   blk00000181 (
    .CI(sig00000283),
    .LI(sig000002fa),
    .O(sig000002c4)
  );
  MUXCY   blk00000182 (
    .CI(sig00000284),
    .DI(sig00000192),
    .S(sig000002fb),
    .O(sig00000285)
  );
  XORCY   blk00000183 (
    .CI(sig00000284),
    .LI(sig000002fb),
    .O(sig000002c5)
  );
  MUXCY   blk00000184 (
    .CI(sig00000285),
    .DI(sig00000193),
    .S(sig000002fc),
    .O(sig00000286)
  );
  XORCY   blk00000185 (
    .CI(sig00000285),
    .LI(sig000002fc),
    .O(sig000002c6)
  );
  MUXCY   blk00000186 (
    .CI(sig00000286),
    .DI(sig00000194),
    .S(sig000002fd),
    .O(sig00000287)
  );
  XORCY   blk00000187 (
    .CI(sig00000286),
    .LI(sig000002fd),
    .O(sig000002c7)
  );
  MUXCY   blk00000188 (
    .CI(sig00000287),
    .DI(sig00000195),
    .S(sig000002fe),
    .O(sig00000288)
  );
  XORCY   blk00000189 (
    .CI(sig00000287),
    .LI(sig000002fe),
    .O(sig000002c8)
  );
  MUXCY   blk0000018a (
    .CI(sig00000288),
    .DI(sig00000196),
    .S(sig000002ff),
    .O(sig00000289)
  );
  XORCY   blk0000018b (
    .CI(sig00000288),
    .LI(sig000002ff),
    .O(sig000002c9)
  );
  MUXCY   blk0000018c (
    .CI(sig00000289),
    .DI(sig00000197),
    .S(sig00000300),
    .O(sig0000028a)
  );
  XORCY   blk0000018d (
    .CI(sig00000289),
    .LI(sig00000300),
    .O(sig000002ca)
  );
  MUXCY   blk0000018e (
    .CI(sig0000028a),
    .DI(sig00000198),
    .S(sig00000301),
    .O(sig0000028b)
  );
  XORCY   blk0000018f (
    .CI(sig0000028a),
    .LI(sig00000301),
    .O(sig000002cb)
  );
  MUXCY   blk00000190 (
    .CI(sig0000028b),
    .DI(sig00000199),
    .S(sig00000302),
    .O(sig0000028c)
  );
  XORCY   blk00000191 (
    .CI(sig0000028b),
    .LI(sig00000302),
    .O(sig000002cc)
  );
  MUXCY   blk00000192 (
    .CI(sig0000028c),
    .DI(sig0000019a),
    .S(sig00000303),
    .O(sig0000028e)
  );
  XORCY   blk00000193 (
    .CI(sig0000028c),
    .LI(sig00000303),
    .O(sig000002cd)
  );
  MUXCY   blk00000194 (
    .CI(sig0000028e),
    .DI(sig0000019c),
    .S(sig00000305),
    .O(sig0000028f)
  );
  XORCY   blk00000195 (
    .CI(sig0000028e),
    .LI(sig00000305),
    .O(sig000002cf)
  );
  MUXCY   blk00000196 (
    .CI(sig0000028f),
    .DI(sig0000019d),
    .S(sig00000306),
    .O(sig00000290)
  );
  XORCY   blk00000197 (
    .CI(sig0000028f),
    .LI(sig00000306),
    .O(sig000002d0)
  );
  MUXCY   blk00000198 (
    .CI(sig00000290),
    .DI(sig0000019e),
    .S(sig00000307),
    .O(sig00000291)
  );
  XORCY   blk00000199 (
    .CI(sig00000290),
    .LI(sig00000307),
    .O(sig000002d1)
  );
  MUXCY   blk0000019a (
    .CI(sig00000291),
    .DI(sig0000019f),
    .S(sig00000308),
    .O(sig00000292)
  );
  XORCY   blk0000019b (
    .CI(sig00000291),
    .LI(sig00000308),
    .O(sig000002d2)
  );
  MUXCY   blk0000019c (
    .CI(sig00000292),
    .DI(sig000001a0),
    .S(sig00000309),
    .O(sig00000293)
  );
  XORCY   blk0000019d (
    .CI(sig00000292),
    .LI(sig00000309),
    .O(sig000002d3)
  );
  MUXCY   blk0000019e (
    .CI(sig00000293),
    .DI(sig000001a1),
    .S(sig0000030a),
    .O(sig00000294)
  );
  XORCY   blk0000019f (
    .CI(sig00000293),
    .LI(sig0000030a),
    .O(sig000002d4)
  );
  MUXCY   blk000001a0 (
    .CI(sig00000294),
    .DI(sig000001a2),
    .S(sig0000030b),
    .O(sig00000295)
  );
  XORCY   blk000001a1 (
    .CI(sig00000294),
    .LI(sig0000030b),
    .O(sig000002d5)
  );
  MUXCY   blk000001a2 (
    .CI(sig00000295),
    .DI(sig000001a3),
    .S(sig0000030c),
    .O(sig00000296)
  );
  XORCY   blk000001a3 (
    .CI(sig00000295),
    .LI(sig0000030c),
    .O(sig000002d6)
  );
  XORCY   blk000001a4 (
    .CI(sig00000296),
    .LI(sig00000280),
    .O(sig000002d7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a5 (
    .C(clk),
    .D(sig000002c3),
    .Q(sig000002a0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a6 (
    .C(clk),
    .D(sig000002ce),
    .Q(sig000002a1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a7 (
    .C(clk),
    .D(sig000002d8),
    .Q(sig000002ac)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a8 (
    .C(clk),
    .D(sig000002d9),
    .Q(sig000002b6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a9 (
    .C(clk),
    .D(sig000002da),
    .Q(sig000002b7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001aa (
    .C(clk),
    .D(sig000002db),
    .Q(sig000002b8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ab (
    .C(clk),
    .D(sig000002dc),
    .Q(sig000002b9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ac (
    .C(clk),
    .D(sig000002dd),
    .Q(sig000002ba)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ad (
    .C(clk),
    .D(sig000002de),
    .Q(sig000002bb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ae (
    .C(clk),
    .D(sig000002df),
    .Q(sig000002bc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001af (
    .C(clk),
    .D(sig000002c4),
    .Q(sig000002a2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b0 (
    .C(clk),
    .D(sig000002c5),
    .Q(sig000002a3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b1 (
    .C(clk),
    .D(sig000002c6),
    .Q(sig000002a4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b2 (
    .C(clk),
    .D(sig000002c7),
    .Q(sig000002a5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b3 (
    .C(clk),
    .D(sig000002c8),
    .Q(sig000002a6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b4 (
    .C(clk),
    .D(sig000002c9),
    .Q(sig000002a7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b5 (
    .C(clk),
    .D(sig000002ca),
    .Q(sig000002a8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b6 (
    .C(clk),
    .D(sig000002cb),
    .Q(sig000002a9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b7 (
    .C(clk),
    .D(sig000002cc),
    .Q(sig000002aa)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b8 (
    .C(clk),
    .D(sig000002cd),
    .Q(sig000002ab)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b9 (
    .C(clk),
    .D(sig000002cf),
    .Q(sig000002ad)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ba (
    .C(clk),
    .D(sig000002d0),
    .Q(sig000002ae)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001bb (
    .C(clk),
    .D(sig000002d1),
    .Q(sig000002af)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001bc (
    .C(clk),
    .D(sig000002d2),
    .Q(sig000002b0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001bd (
    .C(clk),
    .D(sig000002d3),
    .Q(sig000002b1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001be (
    .C(clk),
    .D(sig000002d4),
    .Q(sig000002b2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001bf (
    .C(clk),
    .D(sig000002d5),
    .Q(sig000002b3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c0 (
    .C(clk),
    .D(sig000002d6),
    .Q(sig000002b4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c1 (
    .C(clk),
    .D(sig000002d7),
    .Q(sig000002b5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c2 (
    .C(clk),
    .D(sig00000072),
    .Q(sig000001f6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c3 (
    .C(clk),
    .D(sig00000073),
    .Q(sig000001f7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c4 (
    .C(clk),
    .D(sig00000074),
    .Q(sig00000202)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c5 (
    .C(clk),
    .D(sig00000076),
    .Q(sig0000020b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c6 (
    .C(clk),
    .D(sig00000077),
    .Q(sig0000020c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c7 (
    .C(clk),
    .D(sig00000078),
    .Q(sig0000020d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c8 (
    .C(clk),
    .D(sig00000079),
    .Q(sig0000020e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c9 (
    .C(clk),
    .D(sig0000007a),
    .Q(sig0000020f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ca (
    .C(clk),
    .D(sig0000007b),
    .Q(sig00000210)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001cb (
    .C(clk),
    .D(sig0000007c),
    .Q(sig00000211)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001cc (
    .C(clk),
    .D(sig0000007d),
    .Q(sig000001f8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001cd (
    .C(clk),
    .D(sig0000007e),
    .Q(sig000001f9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ce (
    .C(clk),
    .D(sig0000007f),
    .Q(sig000001fa)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001cf (
    .C(clk),
    .D(sig00000081),
    .Q(sig000001fb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d0 (
    .C(clk),
    .D(sig00000082),
    .Q(sig000001fc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d1 (
    .C(clk),
    .D(sig00000083),
    .Q(sig000001fd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d2 (
    .C(clk),
    .D(sig00000084),
    .Q(sig000001fe)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d3 (
    .C(clk),
    .D(sig00000085),
    .Q(sig000001ff)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d4 (
    .C(clk),
    .D(sig00000086),
    .Q(sig00000200)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d5 (
    .C(clk),
    .D(sig00000087),
    .Q(sig00000201)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d6 (
    .C(clk),
    .D(sig00000088),
    .Q(sig00000203)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d7 (
    .C(clk),
    .D(sig00000089),
    .Q(sig00000204)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d8 (
    .C(clk),
    .D(sig0000008a),
    .Q(sig00000205)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d9 (
    .C(clk),
    .D(sig0000008c),
    .Q(sig00000206)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001da (
    .C(clk),
    .D(sig0000008d),
    .Q(sig00000207)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001db (
    .C(clk),
    .D(sig0000008e),
    .Q(sig00000208)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001dc (
    .C(clk),
    .D(sig0000008f),
    .Q(sig00000209)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001dd (
    .C(clk),
    .D(sig00000090),
    .Q(sig0000020a)
  );
  MUXCY   blk000001de (
    .CI(sig000002be),
    .DI(sig00000001),
    .S(sig0000027f),
    .O(sig000002bf)
  );
  MUXCY   blk000001df (
    .CI(sig00000357),
    .DI(sig00000001),
    .S(sig00000002),
    .O(sig000002be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000359),
    .Q(sig00000156)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000357),
    .Q(sig0000029f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000035e),
    .Q(sig000002bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e0),
    .Q(sig00000528)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005ee),
    .Q(sig000005a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e5 (
    .C(clk),
    .CE(sig00000002),
    .D(b[63]),
    .Q(sig0000046c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e6 (
    .C(clk),
    .CE(sig00000002),
    .D(a[63]),
    .Q(sig00000454)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005eb),
    .Q(sig000005a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005d7),
    .Q(sig0000051b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005d6),
    .Q(sig0000051c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ea (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005ea),
    .Q(sig000004da)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001eb (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005a5),
    .Q(sig000004d5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ec (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005a8),
    .Q(sig000004d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ed (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005aa),
    .Q(sig000004d6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ee (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005a7),
    .Q(sig000004d2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ef (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005a4),
    .Q(sig000004d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005a9),
    .Q(sig000004d4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000008bb),
    .Q(sig000004d1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000046e),
    .Q(sig0000046d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000627),
    .Q(sig0000046e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001f4 (
    .C(clk),
    .D(sig000005db),
    .Q(sig000004ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000049a),
    .Q(sig00000486)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000499),
    .Q(sig00000485)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000484),
    .Q(sig00000470)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000483),
    .Q(sig0000046f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000001f9 (
    .I0(b[52]),
    .I1(a[52]),
    .O(sig000004f8)
  );
  MUXCY   blk000001fa (
    .CI(sig00000002),
    .DI(b[52]),
    .S(sig000004f8),
    .O(sig000004ed)
  );
  XORCY   blk000001fb (
    .CI(sig00000002),
    .LI(sig000004f8),
    .O(sig000005ad)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000001fc (
    .I0(b[53]),
    .I1(a[53]),
    .O(sig000004fa)
  );
  MUXCY   blk000001fd (
    .CI(sig000004ed),
    .DI(b[53]),
    .S(sig000004fa),
    .O(sig000004ef)
  );
  XORCY   blk000001fe (
    .CI(sig000004ed),
    .LI(sig000004fa),
    .O(sig000005b0)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000001ff (
    .I0(b[54]),
    .I1(a[54]),
    .O(sig000004fb)
  );
  MUXCY   blk00000200 (
    .CI(sig000004ef),
    .DI(b[54]),
    .S(sig000004fb),
    .O(sig000004f0)
  );
  XORCY   blk00000201 (
    .CI(sig000004ef),
    .LI(sig000004fb),
    .O(sig000005b1)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000202 (
    .I0(b[55]),
    .I1(a[55]),
    .O(sig000004fc)
  );
  MUXCY   blk00000203 (
    .CI(sig000004f0),
    .DI(b[55]),
    .S(sig000004fc),
    .O(sig000004f1)
  );
  XORCY   blk00000204 (
    .CI(sig000004f0),
    .LI(sig000004fc),
    .O(sig000005b2)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000205 (
    .I0(b[56]),
    .I1(a[56]),
    .O(sig000004fd)
  );
  MUXCY   blk00000206 (
    .CI(sig000004f1),
    .DI(b[56]),
    .S(sig000004fd),
    .O(sig000004f2)
  );
  XORCY   blk00000207 (
    .CI(sig000004f1),
    .LI(sig000004fd),
    .O(sig000005b3)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000208 (
    .I0(b[57]),
    .I1(a[57]),
    .O(sig000004fe)
  );
  MUXCY   blk00000209 (
    .CI(sig000004f2),
    .DI(b[57]),
    .S(sig000004fe),
    .O(sig000004f3)
  );
  XORCY   blk0000020a (
    .CI(sig000004f2),
    .LI(sig000004fe),
    .O(sig000005b4)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000020b (
    .I0(b[58]),
    .I1(a[58]),
    .O(sig000004ff)
  );
  MUXCY   blk0000020c (
    .CI(sig000004f3),
    .DI(b[58]),
    .S(sig000004ff),
    .O(sig000004f4)
  );
  XORCY   blk0000020d (
    .CI(sig000004f3),
    .LI(sig000004ff),
    .O(sig000005b5)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000020e (
    .I0(b[59]),
    .I1(a[59]),
    .O(sig00000500)
  );
  MUXCY   blk0000020f (
    .CI(sig000004f4),
    .DI(b[59]),
    .S(sig00000500),
    .O(sig000004f5)
  );
  XORCY   blk00000210 (
    .CI(sig000004f4),
    .LI(sig00000500),
    .O(sig000005b6)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000211 (
    .I0(b[60]),
    .I1(a[60]),
    .O(sig00000501)
  );
  MUXCY   blk00000212 (
    .CI(sig000004f5),
    .DI(b[60]),
    .S(sig00000501),
    .O(sig000004f6)
  );
  XORCY   blk00000213 (
    .CI(sig000004f5),
    .LI(sig00000501),
    .O(sig000005b7)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000214 (
    .I0(b[61]),
    .I1(a[61]),
    .O(sig00000502)
  );
  MUXCY   blk00000215 (
    .CI(sig000004f6),
    .DI(b[61]),
    .S(sig00000502),
    .O(sig000004f7)
  );
  XORCY   blk00000216 (
    .CI(sig000004f6),
    .LI(sig00000502),
    .O(sig000005b8)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000217 (
    .I0(b[62]),
    .I1(a[62]),
    .O(sig000004f9)
  );
  MUXCY   blk00000218 (
    .CI(sig000004f7),
    .DI(b[62]),
    .S(sig000004f9),
    .O(sig000004ee)
  );
  XORCY   blk00000219 (
    .CI(sig000004f7),
    .LI(sig000004f9),
    .O(sig000005ae)
  );
  XORCY   blk0000021a (
    .CI(sig000004ee),
    .LI(sig00000002),
    .O(sig000005af)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000021b (
    .I0(sig000004c2),
    .I1(sig0000065d),
    .O(sig0000050e)
  );
  MUXCY   blk0000021c (
    .CI(sig00000002),
    .DI(sig000004c2),
    .S(sig0000050e),
    .O(sig00000503)
  );
  XORCY   blk0000021d (
    .CI(sig00000002),
    .LI(sig0000050e),
    .O(sig000005de)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000021e (
    .I0(sig000004c3),
    .I1(sig0000065e),
    .O(sig00000510)
  );
  MUXCY   blk0000021f (
    .CI(sig00000503),
    .DI(sig000004c3),
    .S(sig00000510),
    .O(sig00000505)
  );
  XORCY   blk00000220 (
    .CI(sig00000503),
    .LI(sig00000510),
    .O(sig000005e1)
  );
  MUXCY   blk00000221 (
    .CI(sig00000505),
    .DI(sig000004c5),
    .S(sig00000511),
    .O(sig00000506)
  );
  XORCY   blk00000222 (
    .CI(sig00000505),
    .LI(sig00000511),
    .O(sig000005e2)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000223 (
    .I0(sig000004c6),
    .I1(sig0000065b),
    .O(sig00000512)
  );
  MUXCY   blk00000224 (
    .CI(sig00000506),
    .DI(sig000004c6),
    .S(sig00000512),
    .O(sig00000507)
  );
  XORCY   blk00000225 (
    .CI(sig00000506),
    .LI(sig00000512),
    .O(sig000005e3)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000226 (
    .I0(sig000004c7),
    .I1(sig0000062b),
    .O(sig00000513)
  );
  MUXCY   blk00000227 (
    .CI(sig00000507),
    .DI(sig000004c7),
    .S(sig00000513),
    .O(sig00000508)
  );
  XORCY   blk00000228 (
    .CI(sig00000507),
    .LI(sig00000513),
    .O(sig000005e4)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000229 (
    .I0(sig000004c8),
    .I1(sig0000062a),
    .O(sig00000514)
  );
  MUXCY   blk0000022a (
    .CI(sig00000508),
    .DI(sig000004c8),
    .S(sig00000514),
    .O(sig00000509)
  );
  XORCY   blk0000022b (
    .CI(sig00000508),
    .LI(sig00000514),
    .O(sig000005e5)
  );
  MUXCY   blk0000022c (
    .CI(sig00000509),
    .DI(sig000004c9),
    .S(sig00000515),
    .O(sig0000050a)
  );
  XORCY   blk0000022d (
    .CI(sig00000509),
    .LI(sig00000515),
    .O(sig000005e6)
  );
  MUXCY   blk0000022e (
    .CI(sig0000050a),
    .DI(sig000004ca),
    .S(sig00000516),
    .O(sig0000050b)
  );
  XORCY   blk0000022f (
    .CI(sig0000050a),
    .LI(sig00000516),
    .O(sig000005e7)
  );
  MUXCY   blk00000230 (
    .CI(sig0000050b),
    .DI(sig000004cb),
    .S(sig00000517),
    .O(sig0000050c)
  );
  XORCY   blk00000231 (
    .CI(sig0000050b),
    .LI(sig00000517),
    .O(sig000005e8)
  );
  MUXCY   blk00000232 (
    .CI(sig0000050c),
    .DI(sig000004cc),
    .S(sig00000518),
    .O(sig0000050d)
  );
  XORCY   blk00000233 (
    .CI(sig0000050c),
    .LI(sig00000518),
    .O(sig000005e9)
  );
  MUXCY   blk00000234 (
    .CI(sig0000050d),
    .DI(sig000004c4),
    .S(sig0000050f),
    .O(sig00000504)
  );
  XORCY   blk00000235 (
    .CI(sig0000050d),
    .LI(sig0000050f),
    .O(sig000005df)
  );
  XORCY   blk00000236 (
    .CI(sig00000504),
    .LI(sig00000002),
    .O(sig000005e0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000237 (
    .C(clk),
    .D(sig000004ec),
    .Q(sig0000049f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000238 (
    .C(clk),
    .D(sig000005ed),
    .Q(sig0000049e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000239 (
    .C(clk),
    .D(sig000005ba),
    .Q(sig0000049d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000023a (
    .C(clk),
    .D(sig000005b9),
    .Q(sig0000049c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000023b (
    .C(clk),
    .D(sig000005ec),
    .Q(sig0000049b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023c (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000051f),
    .Q(sig000004e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023d (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000527),
    .Q(sig000004eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023e (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000526),
    .Q(sig000004ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023f (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000525),
    .Q(sig000004e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000240 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000524),
    .Q(sig000004e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000241 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000523),
    .Q(sig000004e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000242 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000522),
    .Q(sig000004e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000243 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000521),
    .Q(sig000004e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000244 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000520),
    .Q(sig000004e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000245 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000051e),
    .Q(sig000004e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000246 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000051d),
    .Q(sig000004e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000247 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005df),
    .Q(sig0000051f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000248 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e9),
    .Q(sig00000527)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000249 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e8),
    .Q(sig00000526)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024a (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e7),
    .Q(sig00000525)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024b (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e6),
    .Q(sig00000524)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024c (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e5),
    .Q(sig00000523)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024d (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e4),
    .Q(sig00000522)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024e (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e3),
    .Q(sig00000521)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024f (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e2),
    .Q(sig00000520)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000250 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005e1),
    .Q(sig0000051e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000251 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000005de),
    .Q(sig0000051d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000252 (
    .C(clk),
    .CE(sig00000002),
    .D(b[62]),
    .Q(sig00000463)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000253 (
    .C(clk),
    .CE(sig00000002),
    .D(b[61]),
    .Q(sig0000046b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000254 (
    .C(clk),
    .CE(sig00000002),
    .D(b[60]),
    .Q(sig0000046a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000255 (
    .C(clk),
    .CE(sig00000002),
    .D(b[59]),
    .Q(sig00000469)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000256 (
    .C(clk),
    .CE(sig00000002),
    .D(b[58]),
    .Q(sig00000468)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000257 (
    .C(clk),
    .CE(sig00000002),
    .D(b[57]),
    .Q(sig00000467)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000258 (
    .C(clk),
    .CE(sig00000002),
    .D(b[56]),
    .Q(sig00000466)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000259 (
    .C(clk),
    .CE(sig00000002),
    .D(b[55]),
    .Q(sig00000465)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025a (
    .C(clk),
    .CE(sig00000002),
    .D(b[54]),
    .Q(sig00000464)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025b (
    .C(clk),
    .CE(sig00000002),
    .D(b[53]),
    .Q(sig00000462)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025c (
    .C(clk),
    .CE(sig00000002),
    .D(b[52]),
    .Q(sig00000461)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025d (
    .C(clk),
    .CE(sig00000002),
    .D(a[62]),
    .Q(sig0000044b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025e (
    .C(clk),
    .CE(sig00000002),
    .D(a[61]),
    .Q(sig00000453)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025f (
    .C(clk),
    .CE(sig00000002),
    .D(a[60]),
    .Q(sig00000452)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000260 (
    .C(clk),
    .CE(sig00000002),
    .D(a[59]),
    .Q(sig00000451)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000261 (
    .C(clk),
    .CE(sig00000002),
    .D(a[58]),
    .Q(sig00000450)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000262 (
    .C(clk),
    .CE(sig00000002),
    .D(a[57]),
    .Q(sig0000044f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000263 (
    .C(clk),
    .CE(sig00000002),
    .D(a[56]),
    .Q(sig0000044e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000264 (
    .C(clk),
    .CE(sig00000002),
    .D(a[55]),
    .Q(sig0000044d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000265 (
    .C(clk),
    .CE(sig00000002),
    .D(a[54]),
    .Q(sig0000044c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000266 (
    .C(clk),
    .CE(sig00000002),
    .D(a[53]),
    .Q(sig0000044a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000267 (
    .C(clk),
    .CE(sig00000002),
    .D(a[52]),
    .Q(sig00000449)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000268 (
    .C(clk),
    .D(sig000005af),
    .Q(sig00000458)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000269 (
    .C(clk),
    .D(sig000005ae),
    .Q(sig00000457)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000026a (
    .C(clk),
    .D(sig000005b8),
    .Q(sig00000460)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000026b (
    .C(clk),
    .D(sig000005b7),
    .Q(sig0000045f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000026c (
    .C(clk),
    .D(sig000005b6),
    .Q(sig0000045e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000026d (
    .C(clk),
    .D(sig000005b5),
    .Q(sig0000045d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000026e (
    .C(clk),
    .D(sig000005b4),
    .Q(sig0000045c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000026f (
    .C(clk),
    .D(sig000005b3),
    .Q(sig0000045b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000270 (
    .C(clk),
    .D(sig000005b2),
    .Q(sig0000045a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000271 (
    .C(clk),
    .D(sig000005b1),
    .Q(sig00000459)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000272 (
    .C(clk),
    .D(sig000005b0),
    .Q(sig00000456)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000273 (
    .C(clk),
    .D(sig000005ad),
    .Q(sig00000455)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000274 (
    .C(clk),
    .D(sig000005bb),
    .Q(sig000004d9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000275 (
    .C(clk),
    .D(sig000005c2),
    .Q(sig000004ae)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000276 (
    .C(clk),
    .D(sig000005c1),
    .Q(sig000004ad)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000277 (
    .C(clk),
    .D(sig000005cb),
    .Q(sig000004b6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000278 (
    .C(clk),
    .D(sig000005ca),
    .Q(sig000004b5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000279 (
    .C(clk),
    .D(sig000005c9),
    .Q(sig000004b4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027a (
    .C(clk),
    .D(sig000005c8),
    .Q(sig000004b3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027b (
    .C(clk),
    .D(sig000005c7),
    .Q(sig000004b2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027c (
    .C(clk),
    .D(sig000005c6),
    .Q(sig000004b1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027d (
    .C(clk),
    .D(sig000005c5),
    .Q(sig000004b0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027e (
    .C(clk),
    .D(sig000005c4),
    .Q(sig000004af)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027f (
    .C(clk),
    .D(sig000005c3),
    .Q(sig000004ac)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000280 (
    .C(clk),
    .D(sig000005c0),
    .Q(sig000004ab)
  );
  XORCY   blk00000281 (
    .CI(sig000004a1),
    .LI(sig00000001),
    .O(sig000005c2)
  );
  XORCY   blk00000282 (
    .CI(sig000004a0),
    .LI(sig000005cc),
    .O(sig000005c1)
  );
  MUXCY   blk00000283 (
    .CI(sig000004a0),
    .DI(sig00000001),
    .S(sig000005cc),
    .O(sig000004a1)
  );
  XORCY   blk00000284 (
    .CI(sig000004aa),
    .LI(sig000005d5),
    .O(sig000005cb)
  );
  MUXCY   blk00000285 (
    .CI(sig000004aa),
    .DI(sig00000001),
    .S(sig000005d5),
    .O(sig000004a0)
  );
  XORCY   blk00000286 (
    .CI(sig000004a9),
    .LI(sig000005d4),
    .O(sig000005ca)
  );
  MUXCY   blk00000287 (
    .CI(sig000004a9),
    .DI(sig00000001),
    .S(sig000005d4),
    .O(sig000004aa)
  );
  XORCY   blk00000288 (
    .CI(sig000004a8),
    .LI(sig000005d3),
    .O(sig000005c9)
  );
  MUXCY   blk00000289 (
    .CI(sig000004a8),
    .DI(sig00000001),
    .S(sig000005d3),
    .O(sig000004a9)
  );
  XORCY   blk0000028a (
    .CI(sig000004a7),
    .LI(sig000005d2),
    .O(sig000005c8)
  );
  MUXCY   blk0000028b (
    .CI(sig000004a7),
    .DI(sig00000001),
    .S(sig000005d2),
    .O(sig000004a8)
  );
  XORCY   blk0000028c (
    .CI(sig000004a6),
    .LI(sig000005d1),
    .O(sig000005c7)
  );
  MUXCY   blk0000028d (
    .CI(sig000004a6),
    .DI(sig00000001),
    .S(sig000005d1),
    .O(sig000004a7)
  );
  XORCY   blk0000028e (
    .CI(sig000004a5),
    .LI(sig000005d0),
    .O(sig000005c6)
  );
  MUXCY   blk0000028f (
    .CI(sig000004a5),
    .DI(sig00000001),
    .S(sig000005d0),
    .O(sig000004a6)
  );
  XORCY   blk00000290 (
    .CI(sig000004a4),
    .LI(sig000005cf),
    .O(sig000005c5)
  );
  MUXCY   blk00000291 (
    .CI(sig000004a4),
    .DI(sig00000001),
    .S(sig000005cf),
    .O(sig000004a5)
  );
  XORCY   blk00000292 (
    .CI(sig000004a3),
    .LI(sig000005ce),
    .O(sig000005c4)
  );
  MUXCY   blk00000293 (
    .CI(sig000004a3),
    .DI(sig00000001),
    .S(sig000005ce),
    .O(sig000004a4)
  );
  XORCY   blk00000294 (
    .CI(sig000004a2),
    .LI(sig000005cd),
    .O(sig000005c3)
  );
  MUXCY   blk00000295 (
    .CI(sig000004a2),
    .DI(sig00000001),
    .S(sig000005cd),
    .O(sig000004a3)
  );
  XORCY   blk00000296 (
    .CI(sig00000001),
    .LI(sig000005ab),
    .O(sig000005c0)
  );
  MUXCY   blk00000297 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000005ab),
    .O(sig000004a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000298 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000479),
    .Q(sig000005a6)
  );
  MUXCY   blk00000299 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig0000047a),
    .O(sig00000471)
  );
  MUXCY   blk0000029a (
    .CI(sig00000471),
    .DI(sig00000001),
    .S(sig0000047b),
    .O(sig00000472)
  );
  MUXCY   blk0000029b (
    .CI(sig00000472),
    .DI(sig00000001),
    .S(sig0000047c),
    .O(sig00000473)
  );
  MUXCY   blk0000029c (
    .CI(sig00000473),
    .DI(sig00000001),
    .S(sig0000047d),
    .O(sig00000474)
  );
  MUXCY   blk0000029d (
    .CI(sig00000474),
    .DI(sig00000001),
    .S(sig0000047e),
    .O(sig00000475)
  );
  MUXCY   blk0000029e (
    .CI(sig00000475),
    .DI(sig00000001),
    .S(sig0000047f),
    .O(sig00000476)
  );
  MUXCY   blk0000029f (
    .CI(sig00000476),
    .DI(sig00000001),
    .S(sig00000480),
    .O(sig00000477)
  );
  MUXCY   blk000002a0 (
    .CI(sig00000477),
    .DI(sig00000001),
    .S(sig00000481),
    .O(sig00000478)
  );
  MUXCY   blk000002a1 (
    .CI(sig00000478),
    .DI(sig00000001),
    .S(sig00000482),
    .O(sig00000479)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000048f),
    .Q(sig000005ac)
  );
  MUXCY   blk000002a3 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000490),
    .O(sig00000487)
  );
  MUXCY   blk000002a4 (
    .CI(sig00000487),
    .DI(sig00000001),
    .S(sig00000491),
    .O(sig00000488)
  );
  MUXCY   blk000002a5 (
    .CI(sig00000488),
    .DI(sig00000001),
    .S(sig00000492),
    .O(sig00000489)
  );
  MUXCY   blk000002a6 (
    .CI(sig00000489),
    .DI(sig00000001),
    .S(sig00000493),
    .O(sig0000048a)
  );
  MUXCY   blk000002a7 (
    .CI(sig0000048a),
    .DI(sig00000001),
    .S(sig00000494),
    .O(sig0000048b)
  );
  MUXCY   blk000002a8 (
    .CI(sig0000048b),
    .DI(sig00000001),
    .S(sig00000495),
    .O(sig0000048c)
  );
  MUXCY   blk000002a9 (
    .CI(sig0000048c),
    .DI(sig00000001),
    .S(sig00000496),
    .O(sig0000048d)
  );
  MUXCY   blk000002aa (
    .CI(sig0000048d),
    .DI(sig00000001),
    .S(sig00000497),
    .O(sig0000048e)
  );
  MUXCY   blk000002ab (
    .CI(sig0000048e),
    .DI(sig00000001),
    .S(sig00000498),
    .O(sig0000048f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ac (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000052f),
    .Q(sig000005a0)
  );
  MUXCY   blk000002ad (
    .CI(sig00000001),
    .DI(sig00000539),
    .S(sig00000549),
    .O(sig00000530)
  );
  MUXCY   blk000002ae (
    .CI(sig00000530),
    .DI(sig00000540),
    .S(sig00000550),
    .O(sig00000531)
  );
  MUXCY   blk000002af (
    .CI(sig00000531),
    .DI(sig00000541),
    .S(sig00000551),
    .O(sig00000532)
  );
  MUXCY   blk000002b0 (
    .CI(sig00000532),
    .DI(sig00000542),
    .S(sig00000552),
    .O(sig00000533)
  );
  MUXCY   blk000002b1 (
    .CI(sig00000533),
    .DI(sig00000543),
    .S(sig00000553),
    .O(sig00000534)
  );
  MUXCY   blk000002b2 (
    .CI(sig00000534),
    .DI(sig00000544),
    .S(sig00000554),
    .O(sig00000535)
  );
  MUXCY   blk000002b3 (
    .CI(sig00000535),
    .DI(sig00000545),
    .S(sig00000555),
    .O(sig00000536)
  );
  MUXCY   blk000002b4 (
    .CI(sig00000536),
    .DI(sig00000546),
    .S(sig00000556),
    .O(sig00000537)
  );
  MUXCY   blk000002b5 (
    .CI(sig00000537),
    .DI(sig00000547),
    .S(sig00000557),
    .O(sig00000538)
  );
  MUXCY   blk000002b6 (
    .CI(sig00000538),
    .DI(sig00000548),
    .S(sig00000558),
    .O(sig00000529)
  );
  MUXCY   blk000002b7 (
    .CI(sig00000529),
    .DI(sig0000053a),
    .S(sig0000054a),
    .O(sig0000052a)
  );
  MUXCY   blk000002b8 (
    .CI(sig0000052a),
    .DI(sig0000053b),
    .S(sig0000054b),
    .O(sig0000052b)
  );
  MUXCY   blk000002b9 (
    .CI(sig0000052b),
    .DI(sig0000053c),
    .S(sig0000054c),
    .O(sig0000052c)
  );
  MUXCY   blk000002ba (
    .CI(sig0000052c),
    .DI(sig0000053d),
    .S(sig0000054d),
    .O(sig0000052d)
  );
  MUXCY   blk000002bb (
    .CI(sig0000052d),
    .DI(sig0000053e),
    .S(sig0000054e),
    .O(sig0000052e)
  );
  MUXCY   blk000002bc (
    .CI(sig0000052e),
    .DI(sig0000053f),
    .S(sig0000054f),
    .O(sig0000052f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002bd (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000575),
    .Q(sig000005a1)
  );
  MUXCY   blk000002be (
    .CI(sig00000001),
    .DI(sig0000057f),
    .S(sig0000058f),
    .O(sig00000576)
  );
  MUXCY   blk000002bf (
    .CI(sig00000576),
    .DI(sig00000586),
    .S(sig00000596),
    .O(sig00000577)
  );
  MUXCY   blk000002c0 (
    .CI(sig00000577),
    .DI(sig00000587),
    .S(sig00000597),
    .O(sig00000578)
  );
  MUXCY   blk000002c1 (
    .CI(sig00000578),
    .DI(sig00000588),
    .S(sig00000598),
    .O(sig00000579)
  );
  MUXCY   blk000002c2 (
    .CI(sig00000579),
    .DI(sig00000589),
    .S(sig00000599),
    .O(sig0000057a)
  );
  MUXCY   blk000002c3 (
    .CI(sig0000057a),
    .DI(sig0000058a),
    .S(sig0000059a),
    .O(sig0000057b)
  );
  MUXCY   blk000002c4 (
    .CI(sig0000057b),
    .DI(sig0000058b),
    .S(sig0000059b),
    .O(sig0000057c)
  );
  MUXCY   blk000002c5 (
    .CI(sig0000057c),
    .DI(sig0000058c),
    .S(sig0000059c),
    .O(sig0000057d)
  );
  MUXCY   blk000002c6 (
    .CI(sig0000057d),
    .DI(sig0000058d),
    .S(sig0000059d),
    .O(sig0000057e)
  );
  MUXCY   blk000002c7 (
    .CI(sig0000057e),
    .DI(sig0000058e),
    .S(sig0000059e),
    .O(sig0000056f)
  );
  MUXCY   blk000002c8 (
    .CI(sig0000056f),
    .DI(sig00000580),
    .S(sig00000590),
    .O(sig00000570)
  );
  MUXCY   blk000002c9 (
    .CI(sig00000570),
    .DI(sig00000581),
    .S(sig00000591),
    .O(sig00000571)
  );
  MUXCY   blk000002ca (
    .CI(sig00000571),
    .DI(sig00000582),
    .S(sig00000592),
    .O(sig00000572)
  );
  MUXCY   blk000002cb (
    .CI(sig00000572),
    .DI(sig00000583),
    .S(sig00000593),
    .O(sig00000573)
  );
  MUXCY   blk000002cc (
    .CI(sig00000573),
    .DI(sig00000584),
    .S(sig00000594),
    .O(sig00000574)
  );
  MUXCY   blk000002cd (
    .CI(sig00000574),
    .DI(sig00000585),
    .S(sig00000595),
    .O(sig00000575)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ce (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000055a),
    .Q(sig0000059f)
  );
  MUXCY   blk000002cf (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000564),
    .O(sig0000055b)
  );
  MUXCY   blk000002d0 (
    .CI(sig0000055b),
    .DI(sig00000001),
    .S(sig00000566),
    .O(sig0000055c)
  );
  MUXCY   blk000002d1 (
    .CI(sig0000055c),
    .DI(sig00000001),
    .S(sig00000567),
    .O(sig0000055d)
  );
  MUXCY   blk000002d2 (
    .CI(sig0000055d),
    .DI(sig00000001),
    .S(sig00000568),
    .O(sig0000055e)
  );
  MUXCY   blk000002d3 (
    .CI(sig0000055e),
    .DI(sig00000001),
    .S(sig00000569),
    .O(sig0000055f)
  );
  MUXCY   blk000002d4 (
    .CI(sig0000055f),
    .DI(sig00000001),
    .S(sig0000056a),
    .O(sig00000560)
  );
  MUXCY   blk000002d5 (
    .CI(sig00000560),
    .DI(sig00000001),
    .S(sig0000056b),
    .O(sig00000561)
  );
  MUXCY   blk000002d6 (
    .CI(sig00000561),
    .DI(sig00000001),
    .S(sig0000056c),
    .O(sig00000562)
  );
  MUXCY   blk000002d7 (
    .CI(sig00000562),
    .DI(sig00000001),
    .S(sig0000056d),
    .O(sig00000563)
  );
  MUXCY   blk000002d8 (
    .CI(sig00000563),
    .DI(sig00000001),
    .S(sig0000056e),
    .O(sig00000559)
  );
  MUXCY   blk000002d9 (
    .CI(sig00000559),
    .DI(sig00000001),
    .S(sig00000565),
    .O(sig0000055a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002da (
    .C(clk),
    .D(sig0000065e),
    .Q(sig00000852)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002db (
    .C(clk),
    .D(sig0000065d),
    .Q(sig00000851)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002dc (
    .C(clk),
    .D(sig000006c8),
    .Q(sig00000849)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002dd (
    .C(clk),
    .D(sig000006d3),
    .Q(sig00000848)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002de (
    .C(clk),
    .D(sig000006de),
    .Q(sig00000847)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002df (
    .C(clk),
    .D(sig000006e9),
    .Q(sig00000846)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e0 (
    .C(clk),
    .D(sig000006f4),
    .Q(sig00000845)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e1 (
    .C(clk),
    .D(sig000006fb),
    .Q(sig00000844)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e2 (
    .C(clk),
    .D(sig000006fc),
    .Q(sig00000843)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e3 (
    .C(clk),
    .D(sig000006fd),
    .Q(sig00000842)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e4 (
    .C(clk),
    .D(sig000006fe),
    .Q(sig00000841)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e5 (
    .C(clk),
    .D(sig000006c9),
    .Q(sig0000083f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e6 (
    .C(clk),
    .D(sig000006ca),
    .Q(sig0000083e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e7 (
    .C(clk),
    .D(sig000006cb),
    .Q(sig0000083d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e8 (
    .C(clk),
    .D(sig000006cc),
    .Q(sig0000083c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002e9 (
    .C(clk),
    .D(sig000006cd),
    .Q(sig0000083b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ea (
    .C(clk),
    .D(sig000006ce),
    .Q(sig0000083a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002eb (
    .C(clk),
    .D(sig000006cf),
    .Q(sig00000839)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ec (
    .C(clk),
    .D(sig000006d0),
    .Q(sig00000838)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ed (
    .C(clk),
    .D(sig000006d1),
    .Q(sig00000837)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ee (
    .C(clk),
    .D(sig000006d2),
    .Q(sig00000836)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ef (
    .C(clk),
    .D(sig000006d4),
    .Q(sig00000850)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f0 (
    .C(clk),
    .D(sig000006d5),
    .Q(sig0000084f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f1 (
    .C(clk),
    .D(sig000006d6),
    .Q(sig0000084e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f2 (
    .C(clk),
    .D(sig000006d7),
    .Q(sig0000084d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f3 (
    .C(clk),
    .D(sig000006d8),
    .Q(sig0000084c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f4 (
    .C(clk),
    .D(sig000006d9),
    .Q(sig0000084b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f5 (
    .C(clk),
    .D(sig000006da),
    .Q(sig0000084a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f6 (
    .C(clk),
    .D(sig000006db),
    .Q(sig00000840)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f7 (
    .C(clk),
    .D(sig000006dc),
    .Q(sig00000835)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002f8 (
    .C(clk),
    .D(sig000006dd),
    .Q(sig00000834)
  );
  XORCY   blk000002f9 (
    .CI(sig0000076d),
    .LI(sig00000001),
    .O(NLW_blk000002f9_O_UNCONNECTED)
  );
  XORCY   blk000002fa (
    .CI(sig00000776),
    .LI(sig00000001),
    .O(NLW_blk000002fa_O_UNCONNECTED)
  );
  MUXCY   blk000002fb (
    .CI(sig00000776),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig0000076d)
  );
  XORCY   blk000002fc (
    .CI(sig00000775),
    .LI(sig00000001),
    .O(NLW_blk000002fc_O_UNCONNECTED)
  );
  MUXCY   blk000002fd (
    .CI(sig00000775),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig00000776)
  );
  XORCY   blk000002fe (
    .CI(sig00000774),
    .LI(sig00000001),
    .O(NLW_blk000002fe_O_UNCONNECTED)
  );
  MUXCY   blk000002ff (
    .CI(sig00000774),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig00000775)
  );
  XORCY   blk00000300 (
    .CI(sig00000773),
    .LI(sig00000001),
    .O(NLW_blk00000300_O_UNCONNECTED)
  );
  MUXCY   blk00000301 (
    .CI(sig00000773),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig00000774)
  );
  XORCY   blk00000302 (
    .CI(sig00000772),
    .LI(sig00000001),
    .O(NLW_blk00000302_O_UNCONNECTED)
  );
  MUXCY   blk00000303 (
    .CI(sig00000772),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig00000773)
  );
  XORCY   blk00000304 (
    .CI(sig00000771),
    .LI(sig00000001),
    .O(NLW_blk00000304_O_UNCONNECTED)
  );
  MUXCY   blk00000305 (
    .CI(sig00000771),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig00000772)
  );
  XORCY   blk00000306 (
    .CI(sig00000770),
    .LI(sig00000001),
    .O(NLW_blk00000306_O_UNCONNECTED)
  );
  MUXCY   blk00000307 (
    .CI(sig00000770),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig00000771)
  );
  XORCY   blk00000308 (
    .CI(sig0000076f),
    .LI(sig00000001),
    .O(NLW_blk00000308_O_UNCONNECTED)
  );
  MUXCY   blk00000309 (
    .CI(sig0000076f),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig00000770)
  );
  XORCY   blk0000030a (
    .CI(sig0000076e),
    .LI(sig00000001),
    .O(NLW_blk0000030a_O_UNCONNECTED)
  );
  MUXCY   blk0000030b (
    .CI(sig0000076e),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig0000076f)
  );
  XORCY   blk0000030c (
    .CI(sig0000085c),
    .LI(sig00000001),
    .O(NLW_blk0000030c_O_UNCONNECTED)
  );
  MUXCY   blk0000030d (
    .CI(sig0000085c),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig0000076e)
  );
  MUXCY   blk0000030e (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000859),
    .O(sig00000854)
  );
  MUXCY   blk0000030f (
    .CI(sig00000854),
    .DI(sig00000002),
    .S(sig0000085a),
    .O(sig00000855)
  );
  MUXCY   blk00000310 (
    .CI(sig00000855),
    .DI(sig00000002),
    .S(sig00000853),
    .O(sig00000856)
  );
  MUXCY   blk00000311 (
    .CI(sig00000856),
    .DI(sig00000001),
    .S(sig0000085b),
    .O(sig00000857)
  );
  MUXCY   blk00000312 (
    .CI(sig00000857),
    .DI(sig00000001),
    .S(sig00000002),
    .O(sig00000858)
  );
  MUXCY   blk00000313 (
    .CI(sig00000858),
    .DI(sig00000002),
    .S(sig00000002),
    .O(sig00000892)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000314 (
    .C(clk),
    .D(sig000007c6),
    .Q(sig00000791)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000315 (
    .C(clk),
    .D(sig000007d1),
    .Q(sig00000792)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000316 (
    .C(clk),
    .D(sig000007d8),
    .Q(sig0000079d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000317 (
    .C(clk),
    .D(sig000007d9),
    .Q(sig000007a4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000318 (
    .C(clk),
    .D(sig000007da),
    .Q(sig000007a5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000319 (
    .C(clk),
    .D(sig000007db),
    .Q(sig000007a6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000031a (
    .C(clk),
    .D(sig000007dc),
    .Q(sig000007a7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000031b (
    .C(clk),
    .D(sig000007dd),
    .Q(sig000007a8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000031c (
    .C(clk),
    .D(sig000007de),
    .Q(sig000007a9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000031d (
    .C(clk),
    .D(sig000007df),
    .Q(sig000007aa)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000031e (
    .C(clk),
    .D(sig000007c7),
    .Q(sig00000793)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000031f (
    .C(clk),
    .D(sig000007c8),
    .Q(sig00000794)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000320 (
    .C(clk),
    .D(sig000007c9),
    .Q(sig00000795)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000321 (
    .C(clk),
    .D(sig000007ca),
    .Q(sig00000796)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000322 (
    .C(clk),
    .D(sig000007cb),
    .Q(sig00000797)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000323 (
    .C(clk),
    .D(sig000007cc),
    .Q(sig00000798)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000324 (
    .C(clk),
    .D(sig000007cd),
    .Q(sig00000799)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000325 (
    .C(clk),
    .D(sig000007ce),
    .Q(sig0000079a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000326 (
    .C(clk),
    .D(sig000007cf),
    .Q(sig0000079b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000327 (
    .C(clk),
    .D(sig000007d0),
    .Q(sig0000079c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000328 (
    .C(clk),
    .D(sig000007d2),
    .Q(sig0000079e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000329 (
    .C(clk),
    .D(sig000007d3),
    .Q(sig0000079f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000032a (
    .C(clk),
    .D(sig000007d4),
    .Q(sig000007a0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000032b (
    .C(clk),
    .D(sig000007d5),
    .Q(sig000007a1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000032c (
    .C(clk),
    .D(sig000007d6),
    .Q(sig000007a2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000032d (
    .C(clk),
    .D(sig000007d7),
    .Q(sig000007a3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000032e (
    .C(clk),
    .D(sig00000791),
    .Q(sig00000777)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000032f (
    .C(clk),
    .D(sig00000792),
    .Q(sig00000778)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000330 (
    .C(clk),
    .D(sig0000079d),
    .Q(sig00000783)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000331 (
    .C(clk),
    .D(sig000007a4),
    .Q(sig0000078a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000332 (
    .C(clk),
    .D(sig000007a5),
    .Q(sig0000078b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000333 (
    .C(clk),
    .D(sig000007a6),
    .Q(sig0000078c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000334 (
    .C(clk),
    .D(sig000007a7),
    .Q(sig0000078d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000335 (
    .C(clk),
    .D(sig000007a8),
    .Q(sig0000078e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000336 (
    .C(clk),
    .D(sig000007a9),
    .Q(sig0000078f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000337 (
    .C(clk),
    .D(sig000007aa),
    .Q(sig00000790)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000338 (
    .C(clk),
    .D(sig00000793),
    .Q(sig00000779)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000339 (
    .C(clk),
    .D(sig00000794),
    .Q(sig0000077a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000033a (
    .C(clk),
    .D(sig00000795),
    .Q(sig0000077b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000033b (
    .C(clk),
    .D(sig00000796),
    .Q(sig0000077c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000033c (
    .C(clk),
    .D(sig00000797),
    .Q(sig0000077d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000033d (
    .C(clk),
    .D(sig00000798),
    .Q(sig0000077e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000033e (
    .C(clk),
    .D(sig00000799),
    .Q(sig0000077f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000033f (
    .C(clk),
    .D(sig0000079a),
    .Q(sig00000780)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000340 (
    .C(clk),
    .D(sig0000079b),
    .Q(sig00000781)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000341 (
    .C(clk),
    .D(sig0000079c),
    .Q(sig00000782)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000342 (
    .C(clk),
    .D(sig0000079e),
    .Q(sig00000784)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000343 (
    .C(clk),
    .D(sig0000079f),
    .Q(sig00000785)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000344 (
    .C(clk),
    .D(sig000007a0),
    .Q(sig00000786)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000345 (
    .C(clk),
    .D(sig000007a1),
    .Q(sig00000787)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000346 (
    .C(clk),
    .D(sig000007a2),
    .Q(sig00000788)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000347 (
    .C(clk),
    .D(sig000007a3),
    .Q(sig00000789)
  );
  XORCY   blk00000348 (
    .CI(sig000007bc),
    .LI(sig00000001),
    .O(sig000007c5)
  );
  XORCY   blk00000349 (
    .CI(sig000007bb),
    .LI(sig0000086f),
    .O(sig000007d7)
  );
  MUXCY   blk0000034a (
    .CI(sig000007bb),
    .DI(sig00000001),
    .S(sig0000086f),
    .O(sig000007bc)
  );
  XORCY   blk0000034b (
    .CI(sig000007ba),
    .LI(sig0000086e),
    .O(sig000007d6)
  );
  MUXCY   blk0000034c (
    .CI(sig000007ba),
    .DI(sig00000001),
    .S(sig0000086e),
    .O(sig000007bb)
  );
  XORCY   blk0000034d (
    .CI(sig000007b9),
    .LI(sig0000086d),
    .O(sig000007d5)
  );
  MUXCY   blk0000034e (
    .CI(sig000007b9),
    .DI(sig00000001),
    .S(sig0000086d),
    .O(sig000007ba)
  );
  XORCY   blk0000034f (
    .CI(sig000007b8),
    .LI(sig0000086c),
    .O(sig000007d4)
  );
  MUXCY   blk00000350 (
    .CI(sig000007b8),
    .DI(sig00000001),
    .S(sig0000086c),
    .O(sig000007b9)
  );
  XORCY   blk00000351 (
    .CI(sig000007b7),
    .LI(sig0000086b),
    .O(sig000007d3)
  );
  MUXCY   blk00000352 (
    .CI(sig000007b7),
    .DI(sig00000001),
    .S(sig0000086b),
    .O(sig000007b8)
  );
  XORCY   blk00000353 (
    .CI(sig000007b6),
    .LI(sig0000086a),
    .O(sig000007d2)
  );
  MUXCY   blk00000354 (
    .CI(sig000007b6),
    .DI(sig00000001),
    .S(sig0000086a),
    .O(sig000007b7)
  );
  XORCY   blk00000355 (
    .CI(sig000007b4),
    .LI(sig00000868),
    .O(sig000007d0)
  );
  MUXCY   blk00000356 (
    .CI(sig000007b4),
    .DI(sig00000001),
    .S(sig00000868),
    .O(sig000007b6)
  );
  XORCY   blk00000357 (
    .CI(sig000007b3),
    .LI(sig00000867),
    .O(sig000007cf)
  );
  MUXCY   blk00000358 (
    .CI(sig000007b3),
    .DI(sig00000001),
    .S(sig00000867),
    .O(sig000007b4)
  );
  XORCY   blk00000359 (
    .CI(sig000007b2),
    .LI(sig00000866),
    .O(sig000007ce)
  );
  MUXCY   blk0000035a (
    .CI(sig000007b2),
    .DI(sig00000001),
    .S(sig00000866),
    .O(sig000007b3)
  );
  XORCY   blk0000035b (
    .CI(sig000007b1),
    .LI(sig00000865),
    .O(sig000007cd)
  );
  MUXCY   blk0000035c (
    .CI(sig000007b1),
    .DI(sig00000001),
    .S(sig00000865),
    .O(sig000007b2)
  );
  XORCY   blk0000035d (
    .CI(sig000007b0),
    .LI(sig00000864),
    .O(sig000007cc)
  );
  MUXCY   blk0000035e (
    .CI(sig000007b0),
    .DI(sig00000001),
    .S(sig00000864),
    .O(sig000007b1)
  );
  XORCY   blk0000035f (
    .CI(sig000007af),
    .LI(sig00000863),
    .O(sig000007cb)
  );
  MUXCY   blk00000360 (
    .CI(sig000007af),
    .DI(sig00000001),
    .S(sig00000863),
    .O(sig000007b0)
  );
  XORCY   blk00000361 (
    .CI(sig000007ae),
    .LI(sig00000862),
    .O(sig000007ca)
  );
  MUXCY   blk00000362 (
    .CI(sig000007ae),
    .DI(sig00000001),
    .S(sig00000862),
    .O(sig000007af)
  );
  XORCY   blk00000363 (
    .CI(sig000007ad),
    .LI(sig00000861),
    .O(sig000007c9)
  );
  MUXCY   blk00000364 (
    .CI(sig000007ad),
    .DI(sig00000001),
    .S(sig00000861),
    .O(sig000007ae)
  );
  XORCY   blk00000365 (
    .CI(sig000007ac),
    .LI(sig00000860),
    .O(sig000007c8)
  );
  MUXCY   blk00000366 (
    .CI(sig000007ac),
    .DI(sig00000001),
    .S(sig00000860),
    .O(sig000007ad)
  );
  XORCY   blk00000367 (
    .CI(sig000007ab),
    .LI(sig0000085f),
    .O(sig000007c7)
  );
  MUXCY   blk00000368 (
    .CI(sig000007ab),
    .DI(sig00000001),
    .S(sig0000085f),
    .O(sig000007ac)
  );
  XORCY   blk00000369 (
    .CI(sig000007c4),
    .LI(sig00000877),
    .O(sig000007df)
  );
  MUXCY   blk0000036a (
    .CI(sig000007c4),
    .DI(sig00000001),
    .S(sig00000877),
    .O(sig000007ab)
  );
  XORCY   blk0000036b (
    .CI(sig000007c3),
    .LI(sig00000876),
    .O(sig000007de)
  );
  MUXCY   blk0000036c (
    .CI(sig000007c3),
    .DI(sig00000001),
    .S(sig00000876),
    .O(sig000007c4)
  );
  XORCY   blk0000036d (
    .CI(sig000007c2),
    .LI(sig00000875),
    .O(sig000007dd)
  );
  MUXCY   blk0000036e (
    .CI(sig000007c2),
    .DI(sig00000001),
    .S(sig00000875),
    .O(sig000007c3)
  );
  XORCY   blk0000036f (
    .CI(sig000007c1),
    .LI(sig00000874),
    .O(sig000007dc)
  );
  MUXCY   blk00000370 (
    .CI(sig000007c1),
    .DI(sig00000001),
    .S(sig00000874),
    .O(sig000007c2)
  );
  XORCY   blk00000371 (
    .CI(sig000007c0),
    .LI(sig00000873),
    .O(sig000007db)
  );
  MUXCY   blk00000372 (
    .CI(sig000007c0),
    .DI(sig00000001),
    .S(sig00000873),
    .O(sig000007c1)
  );
  XORCY   blk00000373 (
    .CI(sig000007bf),
    .LI(sig00000872),
    .O(sig000007da)
  );
  MUXCY   blk00000374 (
    .CI(sig000007bf),
    .DI(sig00000001),
    .S(sig00000872),
    .O(sig000007c0)
  );
  XORCY   blk00000375 (
    .CI(sig000007be),
    .LI(sig00000871),
    .O(sig000007d9)
  );
  MUXCY   blk00000376 (
    .CI(sig000007be),
    .DI(sig00000001),
    .S(sig00000871),
    .O(sig000007bf)
  );
  XORCY   blk00000377 (
    .CI(sig000007bd),
    .LI(sig00000870),
    .O(sig000007d8)
  );
  MUXCY   blk00000378 (
    .CI(sig000007bd),
    .DI(sig00000001),
    .S(sig00000870),
    .O(sig000007be)
  );
  XORCY   blk00000379 (
    .CI(sig000007b5),
    .LI(sig00000869),
    .O(sig000007d1)
  );
  MUXCY   blk0000037a (
    .CI(sig000007b5),
    .DI(sig00000001),
    .S(sig00000869),
    .O(sig000007bd)
  );
  XORCY   blk0000037b (
    .CI(sig00000892),
    .LI(sig0000085e),
    .O(sig000007c6)
  );
  MUXCY   blk0000037c (
    .CI(sig00000892),
    .DI(sig00000001),
    .S(sig0000085e),
    .O(sig000007b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037d (
    .C(clk),
    .CE(sig00000002),
    .D(sig000007c5),
    .Q(sig0000085d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000037e (
    .C(clk),
    .D(sig00000819),
    .Q(sig000007e0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000037f (
    .C(clk),
    .D(sig00000824),
    .Q(sig000007e1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000380 (
    .C(clk),
    .D(sig0000082c),
    .Q(sig000007ec)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000381 (
    .C(clk),
    .D(sig0000082d),
    .Q(sig000007f4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000382 (
    .C(clk),
    .D(sig0000082e),
    .Q(sig000007f5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000383 (
    .C(clk),
    .D(sig0000082f),
    .Q(sig000007f6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000384 (
    .C(clk),
    .D(sig00000830),
    .Q(sig000007f7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000385 (
    .C(clk),
    .D(sig00000831),
    .Q(sig000007f8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000386 (
    .C(clk),
    .D(sig00000832),
    .Q(sig000007f9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000387 (
    .C(clk),
    .D(sig00000833),
    .Q(sig000007fa)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000388 (
    .C(clk),
    .D(sig0000081a),
    .Q(sig000007e2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000389 (
    .C(clk),
    .D(sig0000081b),
    .Q(sig000007e3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000038a (
    .C(clk),
    .D(sig0000081c),
    .Q(sig000007e4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000038b (
    .C(clk),
    .D(sig0000081d),
    .Q(sig000007e5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000038c (
    .C(clk),
    .D(sig0000081e),
    .Q(sig000007e6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000038d (
    .C(clk),
    .D(sig0000081f),
    .Q(sig000007e7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000038e (
    .C(clk),
    .D(sig00000820),
    .Q(sig000007e8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000038f (
    .C(clk),
    .D(sig00000821),
    .Q(sig000007e9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000390 (
    .C(clk),
    .D(sig00000822),
    .Q(sig000007ea)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000391 (
    .C(clk),
    .D(sig00000823),
    .Q(sig000007eb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000392 (
    .C(clk),
    .D(sig00000825),
    .Q(sig000007ed)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000393 (
    .C(clk),
    .D(sig00000826),
    .Q(sig000007ee)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000394 (
    .C(clk),
    .D(sig00000827),
    .Q(sig000007ef)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000395 (
    .C(clk),
    .D(sig00000828),
    .Q(sig000007f0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000396 (
    .C(clk),
    .D(sig00000829),
    .Q(sig000007f1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000397 (
    .C(clk),
    .D(sig0000082a),
    .Q(sig000007f2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000398 (
    .C(clk),
    .D(sig0000082b),
    .Q(sig000007f3)
  );
  XORCY   blk00000399 (
    .CI(sig0000080f),
    .LI(sig00000001),
    .O(sig00000818)
  );
  XORCY   blk0000039a (
    .CI(sig0000080e),
    .LI(sig00000002),
    .O(sig0000082b)
  );
  MUXCY   blk0000039b (
    .CI(sig0000080e),
    .DI(sig00000002),
    .S(sig00000002),
    .O(sig0000080f)
  );
  XORCY   blk0000039c (
    .CI(sig0000080d),
    .LI(sig00000889),
    .O(sig0000082a)
  );
  MUXCY   blk0000039d (
    .CI(sig0000080d),
    .DI(sig00000001),
    .S(sig00000889),
    .O(sig0000080e)
  );
  XORCY   blk0000039e (
    .CI(sig0000080c),
    .LI(sig00000888),
    .O(sig00000829)
  );
  MUXCY   blk0000039f (
    .CI(sig0000080c),
    .DI(sig00000001),
    .S(sig00000888),
    .O(sig0000080d)
  );
  XORCY   blk000003a0 (
    .CI(sig0000080b),
    .LI(sig00000887),
    .O(sig00000828)
  );
  MUXCY   blk000003a1 (
    .CI(sig0000080b),
    .DI(sig00000001),
    .S(sig00000887),
    .O(sig0000080c)
  );
  XORCY   blk000003a2 (
    .CI(sig0000080a),
    .LI(sig00000886),
    .O(sig00000827)
  );
  MUXCY   blk000003a3 (
    .CI(sig0000080a),
    .DI(sig00000001),
    .S(sig00000886),
    .O(sig0000080b)
  );
  XORCY   blk000003a4 (
    .CI(sig00000809),
    .LI(sig00000885),
    .O(sig00000826)
  );
  MUXCY   blk000003a5 (
    .CI(sig00000809),
    .DI(sig00000001),
    .S(sig00000885),
    .O(sig0000080a)
  );
  XORCY   blk000003a6 (
    .CI(sig00000808),
    .LI(sig00000884),
    .O(sig00000825)
  );
  MUXCY   blk000003a7 (
    .CI(sig00000808),
    .DI(sig00000001),
    .S(sig00000884),
    .O(sig00000809)
  );
  XORCY   blk000003a8 (
    .CI(sig00000806),
    .LI(sig00000882),
    .O(sig00000823)
  );
  MUXCY   blk000003a9 (
    .CI(sig00000806),
    .DI(sig00000001),
    .S(sig00000882),
    .O(sig00000808)
  );
  XORCY   blk000003aa (
    .CI(sig00000805),
    .LI(sig00000881),
    .O(sig00000822)
  );
  MUXCY   blk000003ab (
    .CI(sig00000805),
    .DI(sig00000001),
    .S(sig00000881),
    .O(sig00000806)
  );
  XORCY   blk000003ac (
    .CI(sig00000804),
    .LI(sig00000880),
    .O(sig00000821)
  );
  MUXCY   blk000003ad (
    .CI(sig00000804),
    .DI(sig00000001),
    .S(sig00000880),
    .O(sig00000805)
  );
  XORCY   blk000003ae (
    .CI(sig00000803),
    .LI(sig0000087f),
    .O(sig00000820)
  );
  MUXCY   blk000003af (
    .CI(sig00000803),
    .DI(sig00000001),
    .S(sig0000087f),
    .O(sig00000804)
  );
  XORCY   blk000003b0 (
    .CI(sig00000802),
    .LI(sig0000087e),
    .O(sig0000081f)
  );
  MUXCY   blk000003b1 (
    .CI(sig00000802),
    .DI(sig00000001),
    .S(sig0000087e),
    .O(sig00000803)
  );
  XORCY   blk000003b2 (
    .CI(sig00000801),
    .LI(sig0000087d),
    .O(sig0000081e)
  );
  MUXCY   blk000003b3 (
    .CI(sig00000801),
    .DI(sig00000001),
    .S(sig0000087d),
    .O(sig00000802)
  );
  XORCY   blk000003b4 (
    .CI(sig00000800),
    .LI(sig0000087c),
    .O(sig0000081d)
  );
  MUXCY   blk000003b5 (
    .CI(sig00000800),
    .DI(sig00000001),
    .S(sig0000087c),
    .O(sig00000801)
  );
  XORCY   blk000003b6 (
    .CI(sig000007ff),
    .LI(sig0000087b),
    .O(sig0000081c)
  );
  MUXCY   blk000003b7 (
    .CI(sig000007ff),
    .DI(sig00000001),
    .S(sig0000087b),
    .O(sig00000800)
  );
  XORCY   blk000003b8 (
    .CI(sig000007fe),
    .LI(sig0000087a),
    .O(sig0000081b)
  );
  MUXCY   blk000003b9 (
    .CI(sig000007fe),
    .DI(sig00000001),
    .S(sig0000087a),
    .O(sig000007ff)
  );
  XORCY   blk000003ba (
    .CI(sig000007fd),
    .LI(sig00000879),
    .O(sig0000081a)
  );
  MUXCY   blk000003bb (
    .CI(sig000007fd),
    .DI(sig00000001),
    .S(sig00000879),
    .O(sig000007fe)
  );
  XORCY   blk000003bc (
    .CI(sig00000817),
    .LI(sig00000891),
    .O(sig00000833)
  );
  MUXCY   blk000003bd (
    .CI(sig00000817),
    .DI(sig00000001),
    .S(sig00000891),
    .O(sig000007fd)
  );
  XORCY   blk000003be (
    .CI(sig00000816),
    .LI(sig00000890),
    .O(sig00000832)
  );
  MUXCY   blk000003bf (
    .CI(sig00000816),
    .DI(sig00000001),
    .S(sig00000890),
    .O(sig00000817)
  );
  XORCY   blk000003c0 (
    .CI(sig00000815),
    .LI(sig0000088f),
    .O(sig00000831)
  );
  MUXCY   blk000003c1 (
    .CI(sig00000815),
    .DI(sig00000001),
    .S(sig0000088f),
    .O(sig00000816)
  );
  XORCY   blk000003c2 (
    .CI(sig00000814),
    .LI(sig0000088e),
    .O(sig00000830)
  );
  MUXCY   blk000003c3 (
    .CI(sig00000814),
    .DI(sig00000001),
    .S(sig0000088e),
    .O(sig00000815)
  );
  XORCY   blk000003c4 (
    .CI(sig00000813),
    .LI(sig0000088d),
    .O(sig0000082f)
  );
  MUXCY   blk000003c5 (
    .CI(sig00000813),
    .DI(sig00000001),
    .S(sig0000088d),
    .O(sig00000814)
  );
  XORCY   blk000003c6 (
    .CI(sig00000812),
    .LI(sig0000088c),
    .O(sig0000082e)
  );
  MUXCY   blk000003c7 (
    .CI(sig00000812),
    .DI(sig00000001),
    .S(sig0000088c),
    .O(sig00000813)
  );
  XORCY   blk000003c8 (
    .CI(sig00000811),
    .LI(sig0000088b),
    .O(sig0000082d)
  );
  MUXCY   blk000003c9 (
    .CI(sig00000811),
    .DI(sig00000001),
    .S(sig0000088b),
    .O(sig00000812)
  );
  XORCY   blk000003ca (
    .CI(sig00000810),
    .LI(sig0000088a),
    .O(sig0000082c)
  );
  MUXCY   blk000003cb (
    .CI(sig00000810),
    .DI(sig00000001),
    .S(sig0000088a),
    .O(sig00000811)
  );
  XORCY   blk000003cc (
    .CI(sig00000807),
    .LI(sig00000883),
    .O(sig00000824)
  );
  MUXCY   blk000003cd (
    .CI(sig00000807),
    .DI(sig00000001),
    .S(sig00000883),
    .O(sig00000810)
  );
  XORCY   blk000003ce (
    .CI(sig000007fc),
    .LI(sig00000878),
    .O(sig00000819)
  );
  MUXCY   blk000003cf (
    .CI(sig000007fc),
    .DI(sig00000001),
    .S(sig00000878),
    .O(sig00000807)
  );
  MUXCY   blk000003d0 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig000007fb),
    .O(sig000007fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000818),
    .Q(sig0000085c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000675),
    .Q(sig00000627)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000895),
    .Q(sig0000065c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000064d),
    .Q(sig0000065b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000663),
    .Q(sig0000065d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000664),
    .Q(sig0000065e)
  );
  MUXF7   blk000003d7 (
    .I0(sig00000660),
    .I1(sig00000662),
    .S(sig0000064d),
    .O(sig00000664)
  );
  MUXF7   blk000003d8 (
    .I0(sig0000065f),
    .I1(sig00000661),
    .S(sig0000064d),
    .O(sig00000663)
  );
  MUXF7   blk000003d9 (
    .I0(sig00000665),
    .I1(sig00000666),
    .S(sig0000064d),
    .O(NLW_blk000003d9_O_UNCONNECTED)
  );
  MUXCY   blk000003da (
    .CI(sig0000066d),
    .DI(sig00000001),
    .S(sig0000068e),
    .O(sig0000066e)
  );
  MUXCY   blk000003db (
    .CI(sig0000066c),
    .DI(sig00000001),
    .S(sig0000068d),
    .O(sig0000066d)
  );
  MUXCY   blk000003dc (
    .CI(sig0000066b),
    .DI(sig00000001),
    .S(sig0000068c),
    .O(sig0000066c)
  );
  MUXCY   blk000003dd (
    .CI(sig0000066a),
    .DI(sig00000001),
    .S(sig0000068b),
    .O(sig0000066b)
  );
  MUXCY   blk000003de (
    .CI(sig00000669),
    .DI(sig00000001),
    .S(sig0000068a),
    .O(sig0000066a)
  );
  MUXCY   blk000003df (
    .CI(sig00000668),
    .DI(sig00000001),
    .S(sig00000689),
    .O(sig00000669)
  );
  MUXCY   blk000003e0 (
    .CI(sig00000667),
    .DI(sig00000001),
    .S(sig00000688),
    .O(sig00000668)
  );
  MUXCY   blk000003e1 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000683),
    .O(sig00000667)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000066e),
    .Q(sig00000897)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000066d),
    .Q(sig00000680)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000066c),
    .Q(sig0000067f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000066b),
    .Q(sig0000067e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000066a),
    .Q(sig0000067d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000669),
    .Q(sig0000067c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000668),
    .Q(sig0000067b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000667),
    .Q(sig00000676)
  );
  MUXCY   blk000003ea (
    .CI(sig00000673),
    .DI(sig00000001),
    .S(sig00000687),
    .O(sig00000674)
  );
  MUXCY   blk000003eb (
    .CI(sig00000672),
    .DI(sig00000001),
    .S(sig00000686),
    .O(sig00000673)
  );
  MUXCY   blk000003ec (
    .CI(sig00000671),
    .DI(sig00000001),
    .S(sig00000685),
    .O(sig00000672)
  );
  MUXCY   blk000003ed (
    .CI(sig00000670),
    .DI(sig00000001),
    .S(sig00000684),
    .O(sig00000671)
  );
  MUXCY   blk000003ee (
    .CI(sig0000066f),
    .DI(sig00000001),
    .S(sig00000690),
    .O(sig00000670)
  );
  MUXCY   blk000003ef (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig0000068f),
    .O(sig0000066f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000674),
    .Q(sig0000067a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000673),
    .Q(sig00000679)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000672),
    .Q(sig00000678)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000671),
    .Q(sig00000677)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000670),
    .Q(sig00000682)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000066f),
    .Q(sig00000681)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f6 (
    .C(clk),
    .D(sig00000644),
    .Q(sig0000062c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f7 (
    .C(clk),
    .D(sig00000645),
    .Q(sig0000062d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f8 (
    .C(clk),
    .D(sig00000646),
    .Q(sig0000062e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f9 (
    .C(clk),
    .D(sig00000647),
    .Q(sig0000062f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003fa (
    .C(clk),
    .D(sig00000648),
    .Q(sig00000630)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003fb (
    .C(clk),
    .D(sig00000649),
    .Q(sig00000631)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003fc (
    .C(clk),
    .D(sig0000064a),
    .Q(sig00000632)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003fd (
    .C(clk),
    .D(sig0000064b),
    .Q(sig00000633)
  );
  MUXF7   blk000003fe (
    .I0(sig0000063b),
    .I1(sig00000643),
    .S(sig00000897),
    .O(sig0000064b)
  );
  MUXF7   blk000003ff (
    .I0(sig0000063a),
    .I1(sig00000642),
    .S(sig00000897),
    .O(sig0000064a)
  );
  MUXF7   blk00000400 (
    .I0(sig00000639),
    .I1(sig00000641),
    .S(sig00000897),
    .O(sig00000649)
  );
  MUXF7   blk00000401 (
    .I0(sig00000638),
    .I1(sig00000640),
    .S(sig00000897),
    .O(sig00000648)
  );
  MUXF7   blk00000402 (
    .I0(sig00000637),
    .I1(sig0000063f),
    .S(sig00000897),
    .O(sig00000647)
  );
  MUXF7   blk00000403 (
    .I0(sig00000636),
    .I1(sig0000063e),
    .S(sig00000897),
    .O(sig00000646)
  );
  MUXF7   blk00000404 (
    .I0(sig00000635),
    .I1(sig0000063d),
    .S(sig00000897),
    .O(sig00000645)
  );
  MUXF7   blk00000405 (
    .I0(sig00000634),
    .I1(sig0000063c),
    .S(sig00000897),
    .O(sig00000644)
  );
  MUXF7   blk00000406 (
    .I0(sig00000653),
    .I1(sig00000001),
    .S(sig00000897),
    .O(sig0000065a)
  );
  MUXF7   blk00000407 (
    .I0(sig00000652),
    .I1(sig00000656),
    .S(sig00000897),
    .O(sig00000659)
  );
  MUXF7   blk00000408 (
    .I0(sig00000651),
    .I1(sig00000655),
    .S(sig00000897),
    .O(sig00000658)
  );
  MUXF7   blk00000409 (
    .I0(sig00000650),
    .I1(sig00000654),
    .S(sig00000897),
    .O(sig00000657)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000040a (
    .C(clk),
    .D(sig00000657),
    .Q(sig0000064c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000040b (
    .C(clk),
    .D(sig00000658),
    .Q(sig0000064d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000040c (
    .C(clk),
    .D(sig00000659),
    .Q(sig0000064e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000040d (
    .C(clk),
    .D(sig0000065a),
    .Q(sig0000064f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000040e (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000730),
    .Q(sig000006fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000040f (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000072f),
    .Q(sig000006f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000410 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000072e),
    .Q(sig000006f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000411 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000072d),
    .Q(sig000006f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000412 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000072c),
    .Q(sig000006f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000413 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000072b),
    .Q(sig000006f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000414 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000729),
    .Q(sig000006f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000415 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000728),
    .Q(sig000006f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000416 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000727),
    .Q(sig000006f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000417 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000726),
    .Q(sig000006f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000418 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000725),
    .Q(sig000006ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000419 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000724),
    .Q(sig000006ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000041a (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000723),
    .Q(sig000006ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000041b (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000722),
    .Q(sig000006ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000041c (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000721),
    .Q(sig000006eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000041d (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000720),
    .Q(sig000006ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000041e (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000071e),
    .Q(sig000006e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000041f (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000071d),
    .Q(sig000006e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000420 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000071c),
    .Q(sig000006e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000421 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000071b),
    .Q(sig000006e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000422 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000071a),
    .Q(sig000006e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000423 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000719),
    .Q(sig000006e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000424 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000718),
    .Q(sig000006e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000425 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000717),
    .Q(sig000006e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000426 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000716),
    .Q(sig000006e0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000427 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000715),
    .Q(sig000006df)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000428 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000713),
    .Q(sig000006dd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000429 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000712),
    .Q(sig000006dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000042a (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000711),
    .Q(sig000006db)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000042b (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000710),
    .Q(sig000006da)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000042c (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000070f),
    .Q(sig000006d9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000042d (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000070e),
    .Q(sig000006d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000042e (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000070d),
    .Q(sig000006d7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000042f (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000070c),
    .Q(sig000006d6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000430 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000070b),
    .Q(sig000006d5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000431 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000070a),
    .Q(sig000006d4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000432 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000708),
    .Q(sig000006d2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000433 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000707),
    .Q(sig000006d1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000434 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000706),
    .Q(sig000006d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000435 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000705),
    .Q(sig000006cf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000436 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000704),
    .Q(sig000006ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000437 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000703),
    .Q(sig000006cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000438 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000702),
    .Q(sig000006cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000439 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000701),
    .Q(sig000006cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000043a (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000700),
    .Q(sig000006ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000043b (
    .C(clk),
    .CE(sig00000002),
    .D(sig000006ff),
    .Q(sig000006c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000043c (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000735),
    .Q(sig000006fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000043d (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000734),
    .Q(sig000006fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000043e (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000733),
    .Q(sig000006fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000043f (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000732),
    .Q(sig000006fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000440 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000731),
    .Q(sig000006f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000441 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000072a),
    .Q(sig000006e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000442 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000071f),
    .Q(sig000006de)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000443 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000714),
    .Q(sig000006d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000444 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000709),
    .Q(sig000006c8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000445 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000767),
    .Q(sig000006c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000446 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000766),
    .Q(sig000006c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000447 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000765),
    .Q(sig000006c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000448 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000764),
    .Q(sig000006c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000449 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000763),
    .Q(sig000006bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000044a (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000762),
    .Q(sig000006be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000044b (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000760),
    .Q(sig000006bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000044c (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000075f),
    .Q(sig000006bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000044d (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000075e),
    .Q(sig000006ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000044e (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000075d),
    .Q(sig000006b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000044f (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000075c),
    .Q(sig000006b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000450 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000075b),
    .Q(sig000006b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000451 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000075a),
    .Q(sig000006b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000452 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000759),
    .Q(sig000006b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000453 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000758),
    .Q(sig000006b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000454 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000757),
    .Q(sig000006b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000455 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000755),
    .Q(sig000006b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000456 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000754),
    .Q(sig000006b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000457 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000753),
    .Q(sig000006af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000458 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000752),
    .Q(sig000006ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000459 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000751),
    .Q(sig000006ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000045a (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000750),
    .Q(sig000006ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000045b (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000074f),
    .Q(sig000006ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000045c (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000074e),
    .Q(sig000006aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000045d (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000074d),
    .Q(sig000006a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000045e (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000074c),
    .Q(sig000006a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000045f (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000074a),
    .Q(sig000006a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000460 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000749),
    .Q(sig000006a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000461 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000748),
    .Q(sig000006a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000462 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000747),
    .Q(sig000006a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000463 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000746),
    .Q(sig000006a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000464 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000745),
    .Q(sig000006a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000465 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000744),
    .Q(sig000006a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000466 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000743),
    .Q(sig0000069f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000467 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000742),
    .Q(sig0000069e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000468 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000741),
    .Q(sig0000069d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000469 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000073f),
    .Q(sig0000069b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000046a (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000073e),
    .Q(sig0000069a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000046b (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000073d),
    .Q(sig00000699)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000046c (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000073c),
    .Q(sig00000698)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000046d (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000073b),
    .Q(sig00000697)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000046e (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000073a),
    .Q(sig00000696)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000046f (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000739),
    .Q(sig00000695)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000470 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000738),
    .Q(sig00000694)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000471 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000737),
    .Q(sig00000693)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000472 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000736),
    .Q(sig00000692)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000473 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000076c),
    .Q(sig000006c7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000474 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000076b),
    .Q(sig000006c6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000475 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000076a),
    .Q(sig000006c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000476 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000769),
    .Q(sig000006c4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000477 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000768),
    .Q(sig000006bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000478 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000761),
    .Q(sig000006b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000479 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000756),
    .Q(sig000006a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000047a (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000074b),
    .Q(sig0000069c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000047b (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000740),
    .Q(sig00000691)
  );
  FDRS   blk0000047c (
    .C(clk),
    .D(sig00000779),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [10])
  );
  FDRS   blk0000047d (
    .C(clk),
    .D(sig0000077a),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [11])
  );
  FDRS   blk0000047e (
    .C(clk),
    .D(sig0000077b),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [12])
  );
  FDRS   blk0000047f (
    .C(clk),
    .D(sig0000077c),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [13])
  );
  FDRS   blk00000480 (
    .C(clk),
    .D(sig0000077d),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [14])
  );
  FDRS   blk00000481 (
    .C(clk),
    .D(sig00000784),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [20])
  );
  FDRS   blk00000482 (
    .C(clk),
    .D(sig0000077e),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [15])
  );
  FDRS   blk00000483 (
    .C(clk),
    .D(sig00000785),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [21])
  );
  FDRS   blk00000484 (
    .C(clk),
    .D(sig0000077f),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [16])
  );
  FDRS   blk00000485 (
    .C(clk),
    .D(sig00000780),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [17])
  );
  FDRS   blk00000486 (
    .C(clk),
    .D(sig00000786),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [22])
  );
  FDRS   blk00000487 (
    .C(clk),
    .D(sig00000787),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [23])
  );
  FDRS   blk00000488 (
    .C(clk),
    .D(sig00000781),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [18])
  );
  FDRS   blk00000489 (
    .C(clk),
    .D(sig00000788),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [24])
  );
  FDRS   blk0000048a (
    .C(clk),
    .D(sig00000782),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [19])
  );
  FDRS   blk0000048b (
    .C(clk),
    .D(sig000007f6),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [31])
  );
  FDRS   blk0000048c (
    .C(clk),
    .D(sig000007f5),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [30])
  );
  FDRS   blk0000048d (
    .C(clk),
    .D(sig00000789),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [25])
  );
  FDRS   blk0000048e (
    .C(clk),
    .D(sig000007e0),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [26])
  );
  FDRS   blk0000048f (
    .C(clk),
    .D(sig00000777),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [0])
  );
  FDRS   blk00000490 (
    .C(clk),
    .D(sig000007f7),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [32])
  );
  FDRS   blk00000491 (
    .C(clk),
    .D(sig000007e1),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [27])
  );
  FDRS   blk00000492 (
    .C(clk),
    .D(sig000007ec),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [28])
  );
  FDRS   blk00000493 (
    .C(clk),
    .D(sig00000778),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [1])
  );
  FDRS   blk00000494 (
    .C(clk),
    .D(sig000007f8),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [33])
  );
  FDRS   blk00000495 (
    .C(clk),
    .D(sig00000783),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [2])
  );
  FDRS   blk00000496 (
    .C(clk),
    .D(sig000007f9),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [34])
  );
  FDRS   blk00000497 (
    .C(clk),
    .D(sig000007f4),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [29])
  );
  FDRS   blk00000498 (
    .C(clk),
    .D(sig0000078a),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [3])
  );
  FDRS   blk00000499 (
    .C(clk),
    .D(sig000007e6),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [40])
  );
  FDRS   blk0000049a (
    .C(clk),
    .D(sig000007fa),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [35])
  );
  FDRS   blk0000049b (
    .C(clk),
    .D(sig0000078b),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [4])
  );
  FDRS   blk0000049c (
    .C(clk),
    .D(sig000007e7),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [41])
  );
  FDRS   blk0000049d (
    .C(clk),
    .D(sig000007e2),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [36])
  );
  FDRS   blk0000049e (
    .C(clk),
    .D(sig0000078c),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [5])
  );
  FDRS   blk0000049f (
    .C(clk),
    .D(sig000007e8),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [42])
  );
  FDRS   blk000004a0 (
    .C(clk),
    .D(sig000007e3),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [37])
  );
  FDRS   blk000004a1 (
    .C(clk),
    .D(sig000007e4),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [38])
  );
  FDRS   blk000004a2 (
    .C(clk),
    .D(sig0000078d),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [6])
  );
  FDRS   blk000004a3 (
    .C(clk),
    .D(sig000007e9),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [43])
  );
  FDRS   blk000004a4 (
    .C(clk),
    .D(sig0000078e),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [7])
  );
  FDRS   blk000004a5 (
    .C(clk),
    .D(sig000007ea),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [44])
  );
  FDRS   blk000004a6 (
    .C(clk),
    .D(sig000007e5),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [39])
  );
  FDRS   blk000004a7 (
    .C(clk),
    .D(sig0000078f),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [8])
  );
  FDRS   blk000004a8 (
    .C(clk),
    .D(sig00000790),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [9])
  );
  FDRS   blk000004a9 (
    .C(clk),
    .D(sig000007f1),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [50])
  );
  FDRS   blk000004aa (
    .C(clk),
    .D(sig000007eb),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [45])
  );
  FDRS   blk000004ab (
    .C(clk),
    .D(sig000007f2),
    .R(sig0000049e),
    .S(sig0000049d),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [51])
  );
  FDRS   blk000004ac (
    .C(clk),
    .D(sig000007ed),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [46])
  );
  FDRS   blk000004ad (
    .C(clk),
    .D(sig000005a2),
    .R(sig00000001),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op )
  );
  FDRS   blk000004ae (
    .C(clk),
    .D(sig000007ee),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [47])
  );
  FDRS   blk000004af (
    .C(clk),
    .D(sig000007ef),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [48])
  );
  FDRS   blk000004b0 (
    .C(clk),
    .D(sig000007f0),
    .R(sig0000049f),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [49])
  );
  FD   blk000004b1 (
    .C(clk),
    .D(sig000008ae),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [0])
  );
  FD   blk000004b2 (
    .C(clk),
    .D(sig000008b0),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [1])
  );
  FD   blk000004b3 (
    .C(clk),
    .D(sig000008b1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [2])
  );
  FD   blk000004b4 (
    .C(clk),
    .D(sig000008b2),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [3])
  );
  FD   blk000004b5 (
    .C(clk),
    .D(sig000008b3),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [4])
  );
  FD   blk000004b6 (
    .C(clk),
    .D(sig000008b4),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [5])
  );
  FD   blk000004b7 (
    .C(clk),
    .D(sig000008b5),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [6])
  );
  FD   blk000004b8 (
    .C(clk),
    .D(sig000008b6),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [7])
  );
  FD   blk000004b9 (
    .C(clk),
    .D(sig000008b7),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [8])
  );
  FD   blk000004ba (
    .C(clk),
    .D(sig000008b8),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [9])
  );
  FD   blk000004bb (
    .C(clk),
    .D(sig000008af),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [10])
  );
  MUXCY   blk000004bc (
    .CI(sig00000001),
    .DI(sig000008a3),
    .S(sig000008a2),
    .O(sig00000898)
  );
  XORCY   blk000004bd (
    .CI(sig00000001),
    .LI(sig000008a2),
    .O(sig000008ae)
  );
  MUXCY   blk000004be (
    .CI(sig00000898),
    .DI(sig00000001),
    .S(sig000008a5),
    .O(sig00000899)
  );
  XORCY   blk000004bf (
    .CI(sig00000898),
    .LI(sig000008a5),
    .O(sig000008b0)
  );
  MUXCY   blk000004c0 (
    .CI(sig00000899),
    .DI(sig00000001),
    .S(sig000008a6),
    .O(sig0000089a)
  );
  XORCY   blk000004c1 (
    .CI(sig00000899),
    .LI(sig000008a6),
    .O(sig000008b1)
  );
  MUXCY   blk000004c2 (
    .CI(sig0000089a),
    .DI(sig00000001),
    .S(sig000008a7),
    .O(sig0000089b)
  );
  XORCY   blk000004c3 (
    .CI(sig0000089a),
    .LI(sig000008a7),
    .O(sig000008b2)
  );
  MUXCY   blk000004c4 (
    .CI(sig0000089b),
    .DI(sig00000001),
    .S(sig000008a8),
    .O(sig0000089c)
  );
  XORCY   blk000004c5 (
    .CI(sig0000089b),
    .LI(sig000008a8),
    .O(sig000008b3)
  );
  MUXCY   blk000004c6 (
    .CI(sig0000089c),
    .DI(sig00000001),
    .S(sig000008a9),
    .O(sig0000089d)
  );
  XORCY   blk000004c7 (
    .CI(sig0000089c),
    .LI(sig000008a9),
    .O(sig000008b4)
  );
  MUXCY   blk000004c8 (
    .CI(sig0000089d),
    .DI(sig00000001),
    .S(sig000008aa),
    .O(sig0000089e)
  );
  XORCY   blk000004c9 (
    .CI(sig0000089d),
    .LI(sig000008aa),
    .O(sig000008b5)
  );
  MUXCY   blk000004ca (
    .CI(sig0000089e),
    .DI(sig00000001),
    .S(sig000008ab),
    .O(sig0000089f)
  );
  XORCY   blk000004cb (
    .CI(sig0000089e),
    .LI(sig000008ab),
    .O(sig000008b6)
  );
  MUXCY   blk000004cc (
    .CI(sig0000089f),
    .DI(sig00000001),
    .S(sig000008ac),
    .O(sig000008a0)
  );
  XORCY   blk000004cd (
    .CI(sig0000089f),
    .LI(sig000008ac),
    .O(sig000008b7)
  );
  MUXCY   blk000004ce (
    .CI(sig000008a0),
    .DI(sig00000001),
    .S(sig000008ad),
    .O(sig000008a1)
  );
  XORCY   blk000004cf (
    .CI(sig000008a0),
    .LI(sig000008ad),
    .O(sig000008b8)
  );
  XORCY   blk000004d0 (
    .CI(sig000008a1),
    .LI(sig000008a4),
    .O(sig000008af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000212),
    .Q(sig000005ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000213),
    .Q(sig000005f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000021e),
    .Q(sig000005fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000226),
    .Q(sig00000606)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000227),
    .Q(sig00000611)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000228),
    .Q(sig0000061c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000229),
    .Q(sig00000623)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000022a),
    .Q(sig00000624)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004d9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000022b),
    .Q(sig00000625)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004da (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000022c),
    .Q(sig00000626)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004db (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000214),
    .Q(sig000005f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004dc (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000215),
    .Q(sig000005f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004dd (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000216),
    .Q(sig000005f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004de (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000217),
    .Q(sig000005f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004df (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000218),
    .Q(sig000005f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000219),
    .Q(sig000005f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000021a),
    .Q(sig000005f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000021b),
    .Q(sig000005f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000021c),
    .Q(sig000005f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000021d),
    .Q(sig000005fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000021f),
    .Q(sig000005fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000220),
    .Q(sig000005fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000221),
    .Q(sig000005fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000222),
    .Q(sig000005ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000223),
    .Q(sig00000600)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ea (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000224),
    .Q(sig00000601)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004eb (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000225),
    .Q(sig00000602)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ec (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a0),
    .Q(sig00000603)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ed (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a1),
    .Q(sig00000604)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ee (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002ac),
    .Q(sig00000605)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ef (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b6),
    .Q(sig00000607)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b7),
    .Q(sig00000608)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f1 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b8),
    .Q(sig00000609)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b9),
    .Q(sig0000060a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f3 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002ba),
    .Q(sig0000060b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002bb),
    .Q(sig0000060c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f5 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002bc),
    .Q(sig0000060d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a2),
    .Q(sig0000060e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f7 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a3),
    .Q(sig0000060f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a4),
    .Q(sig00000610)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f9 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a5),
    .Q(sig00000612)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fa (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a6),
    .Q(sig00000613)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fb (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a7),
    .Q(sig00000614)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fc (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a8),
    .Q(sig00000615)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fd (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002a9),
    .Q(sig00000616)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fe (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002aa),
    .Q(sig00000617)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ff (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002ab),
    .Q(sig00000618)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000500 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002ad),
    .Q(sig00000619)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000501 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002ae),
    .Q(sig0000061a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000502 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002af),
    .Q(sig0000061b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000503 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b0),
    .Q(sig0000061d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000504 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b1),
    .Q(sig0000061e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000505 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b2),
    .Q(sig0000061f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000506 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b3),
    .Q(sig00000620)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000507 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b4),
    .Q(sig00000621)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000508 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000002b5),
    .Q(sig00000622)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000509 (
    .C(clk),
    .CE(sig00000002),
    .D(a[0]),
    .Q(sig000003e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000050a (
    .C(clk),
    .CE(sig00000002),
    .D(a[1]),
    .Q(sig000003e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000050b (
    .C(clk),
    .CE(sig00000002),
    .D(a[2]),
    .Q(sig000003ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000050c (
    .C(clk),
    .CE(sig00000002),
    .D(a[3]),
    .Q(sig000003f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000050d (
    .C(clk),
    .CE(sig00000002),
    .D(a[4]),
    .Q(sig00000403)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000050e (
    .C(clk),
    .CE(sig00000002),
    .D(a[5]),
    .Q(sig0000040e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000050f (
    .C(clk),
    .CE(sig00000002),
    .D(a[6]),
    .Q(sig00000411)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000510 (
    .C(clk),
    .CE(sig00000002),
    .D(a[7]),
    .Q(sig00000412)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000511 (
    .C(clk),
    .CE(sig00000002),
    .D(a[8]),
    .Q(sig00000413)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000512 (
    .C(clk),
    .CE(sig00000002),
    .D(a[9]),
    .Q(sig00000414)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000513 (
    .C(clk),
    .CE(sig00000002),
    .D(a[10]),
    .Q(sig000003e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000514 (
    .C(clk),
    .CE(sig00000002),
    .D(a[11]),
    .Q(sig000003e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000515 (
    .C(clk),
    .CE(sig00000002),
    .D(a[12]),
    .Q(sig000003e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000516 (
    .C(clk),
    .CE(sig00000002),
    .D(a[13]),
    .Q(sig000003e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000517 (
    .C(clk),
    .CE(sig00000002),
    .D(a[14]),
    .Q(sig000003e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000518 (
    .C(clk),
    .CE(sig00000002),
    .D(a[15]),
    .Q(sig000003e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000519 (
    .C(clk),
    .CE(sig00000002),
    .D(a[16]),
    .Q(sig000003e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000051a (
    .C(clk),
    .CE(sig00000002),
    .D(a[17]),
    .Q(sig000003ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000051b (
    .C(clk),
    .CE(sig00000002),
    .D(a[18]),
    .Q(sig000003eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000051c (
    .C(clk),
    .CE(sig00000002),
    .D(a[19]),
    .Q(sig000003ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000051d (
    .C(clk),
    .CE(sig00000002),
    .D(a[20]),
    .Q(sig000003ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000051e (
    .C(clk),
    .CE(sig00000002),
    .D(a[21]),
    .Q(sig000003ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000051f (
    .C(clk),
    .CE(sig00000002),
    .D(a[22]),
    .Q(sig000003f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000520 (
    .C(clk),
    .CE(sig00000002),
    .D(a[23]),
    .Q(sig000003f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000521 (
    .C(clk),
    .CE(sig00000002),
    .D(a[24]),
    .Q(sig000003f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000522 (
    .C(clk),
    .CE(sig00000002),
    .D(a[25]),
    .Q(sig000003f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000523 (
    .C(clk),
    .CE(sig00000002),
    .D(a[26]),
    .Q(sig000003f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000524 (
    .C(clk),
    .CE(sig00000002),
    .D(a[27]),
    .Q(sig000003f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000525 (
    .C(clk),
    .CE(sig00000002),
    .D(a[28]),
    .Q(sig000003f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000526 (
    .C(clk),
    .CE(sig00000002),
    .D(a[29]),
    .Q(sig000003f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000527 (
    .C(clk),
    .CE(sig00000002),
    .D(a[30]),
    .Q(sig000003f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000528 (
    .C(clk),
    .CE(sig00000002),
    .D(a[31]),
    .Q(sig000003fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000529 (
    .C(clk),
    .CE(sig00000002),
    .D(a[32]),
    .Q(sig000003fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000052a (
    .C(clk),
    .CE(sig00000002),
    .D(a[33]),
    .Q(sig000003fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000052b (
    .C(clk),
    .CE(sig00000002),
    .D(a[34]),
    .Q(sig000003fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000052c (
    .C(clk),
    .CE(sig00000002),
    .D(a[35]),
    .Q(sig000003fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000052d (
    .C(clk),
    .CE(sig00000002),
    .D(a[36]),
    .Q(sig000003ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000052e (
    .C(clk),
    .CE(sig00000002),
    .D(a[37]),
    .Q(sig00000400)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000052f (
    .C(clk),
    .CE(sig00000002),
    .D(a[38]),
    .Q(sig00000401)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000530 (
    .C(clk),
    .CE(sig00000002),
    .D(a[39]),
    .Q(sig00000402)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000531 (
    .C(clk),
    .CE(sig00000002),
    .D(a[40]),
    .Q(sig00000404)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000532 (
    .C(clk),
    .CE(sig00000002),
    .D(a[41]),
    .Q(sig00000405)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000533 (
    .C(clk),
    .CE(sig00000002),
    .D(a[42]),
    .Q(sig00000406)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000534 (
    .C(clk),
    .CE(sig00000002),
    .D(a[43]),
    .Q(sig00000407)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000535 (
    .C(clk),
    .CE(sig00000002),
    .D(a[44]),
    .Q(sig00000408)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000536 (
    .C(clk),
    .CE(sig00000002),
    .D(a[45]),
    .Q(sig00000409)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000537 (
    .C(clk),
    .CE(sig00000002),
    .D(a[46]),
    .Q(sig0000040a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000538 (
    .C(clk),
    .CE(sig00000002),
    .D(a[47]),
    .Q(sig0000040b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000539 (
    .C(clk),
    .CE(sig00000002),
    .D(a[48]),
    .Q(sig0000040c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000053a (
    .C(clk),
    .CE(sig00000002),
    .D(a[49]),
    .Q(sig0000040d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000053b (
    .C(clk),
    .CE(sig00000002),
    .D(a[50]),
    .Q(sig0000040f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000053c (
    .C(clk),
    .CE(sig00000002),
    .D(a[51]),
    .Q(sig00000410)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000053d (
    .C(clk),
    .CE(sig00000002),
    .D(b[0]),
    .Q(sig00000415)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000053e (
    .C(clk),
    .CE(sig00000002),
    .D(b[1]),
    .Q(sig00000416)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000053f (
    .C(clk),
    .CE(sig00000002),
    .D(b[2]),
    .Q(sig00000421)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000540 (
    .C(clk),
    .CE(sig00000002),
    .D(b[3]),
    .Q(sig0000042c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000541 (
    .C(clk),
    .CE(sig00000002),
    .D(b[4]),
    .Q(sig00000437)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000542 (
    .C(clk),
    .CE(sig00000002),
    .D(b[5]),
    .Q(sig00000442)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000543 (
    .C(clk),
    .CE(sig00000002),
    .D(b[6]),
    .Q(sig00000445)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000544 (
    .C(clk),
    .CE(sig00000002),
    .D(b[7]),
    .Q(sig00000446)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000545 (
    .C(clk),
    .CE(sig00000002),
    .D(b[8]),
    .Q(sig00000447)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000546 (
    .C(clk),
    .CE(sig00000002),
    .D(b[9]),
    .Q(sig00000448)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000547 (
    .C(clk),
    .CE(sig00000002),
    .D(b[10]),
    .Q(sig00000417)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000548 (
    .C(clk),
    .CE(sig00000002),
    .D(b[11]),
    .Q(sig00000418)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000549 (
    .C(clk),
    .CE(sig00000002),
    .D(b[12]),
    .Q(sig00000419)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000054a (
    .C(clk),
    .CE(sig00000002),
    .D(b[13]),
    .Q(sig0000041a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000054b (
    .C(clk),
    .CE(sig00000002),
    .D(b[14]),
    .Q(sig0000041b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000054c (
    .C(clk),
    .CE(sig00000002),
    .D(b[15]),
    .Q(sig0000041c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000054d (
    .C(clk),
    .CE(sig00000002),
    .D(b[16]),
    .Q(sig0000041d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000054e (
    .C(clk),
    .CE(sig00000002),
    .D(b[17]),
    .Q(sig0000041e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000054f (
    .C(clk),
    .CE(sig00000002),
    .D(b[18]),
    .Q(sig0000041f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000550 (
    .C(clk),
    .CE(sig00000002),
    .D(b[19]),
    .Q(sig00000420)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000551 (
    .C(clk),
    .CE(sig00000002),
    .D(b[20]),
    .Q(sig00000422)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000552 (
    .C(clk),
    .CE(sig00000002),
    .D(b[21]),
    .Q(sig00000423)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000553 (
    .C(clk),
    .CE(sig00000002),
    .D(b[22]),
    .Q(sig00000424)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000554 (
    .C(clk),
    .CE(sig00000002),
    .D(b[23]),
    .Q(sig00000425)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000555 (
    .C(clk),
    .CE(sig00000002),
    .D(b[24]),
    .Q(sig00000426)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000556 (
    .C(clk),
    .CE(sig00000002),
    .D(b[25]),
    .Q(sig00000427)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000557 (
    .C(clk),
    .CE(sig00000002),
    .D(b[26]),
    .Q(sig00000428)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000558 (
    .C(clk),
    .CE(sig00000002),
    .D(b[27]),
    .Q(sig00000429)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000559 (
    .C(clk),
    .CE(sig00000002),
    .D(b[28]),
    .Q(sig0000042a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055a (
    .C(clk),
    .CE(sig00000002),
    .D(b[29]),
    .Q(sig0000042b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055b (
    .C(clk),
    .CE(sig00000002),
    .D(b[30]),
    .Q(sig0000042d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055c (
    .C(clk),
    .CE(sig00000002),
    .D(b[31]),
    .Q(sig0000042e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055d (
    .C(clk),
    .CE(sig00000002),
    .D(b[32]),
    .Q(sig0000042f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055e (
    .C(clk),
    .CE(sig00000002),
    .D(b[33]),
    .Q(sig00000430)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055f (
    .C(clk),
    .CE(sig00000002),
    .D(b[34]),
    .Q(sig00000431)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000560 (
    .C(clk),
    .CE(sig00000002),
    .D(b[35]),
    .Q(sig00000432)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000561 (
    .C(clk),
    .CE(sig00000002),
    .D(b[36]),
    .Q(sig00000433)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000562 (
    .C(clk),
    .CE(sig00000002),
    .D(b[37]),
    .Q(sig00000434)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000563 (
    .C(clk),
    .CE(sig00000002),
    .D(b[38]),
    .Q(sig00000435)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000564 (
    .C(clk),
    .CE(sig00000002),
    .D(b[39]),
    .Q(sig00000436)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000565 (
    .C(clk),
    .CE(sig00000002),
    .D(b[40]),
    .Q(sig00000438)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000566 (
    .C(clk),
    .CE(sig00000002),
    .D(b[41]),
    .Q(sig00000439)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000567 (
    .C(clk),
    .CE(sig00000002),
    .D(b[42]),
    .Q(sig0000043a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000568 (
    .C(clk),
    .CE(sig00000002),
    .D(b[43]),
    .Q(sig0000043b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000569 (
    .C(clk),
    .CE(sig00000002),
    .D(b[44]),
    .Q(sig0000043c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056a (
    .C(clk),
    .CE(sig00000002),
    .D(b[45]),
    .Q(sig0000043d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056b (
    .C(clk),
    .CE(sig00000002),
    .D(b[46]),
    .Q(sig0000043e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056c (
    .C(clk),
    .CE(sig00000002),
    .D(b[47]),
    .Q(sig0000043f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056d (
    .C(clk),
    .CE(sig00000002),
    .D(b[48]),
    .Q(sig00000440)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056e (
    .C(clk),
    .CE(sig00000002),
    .D(b[49]),
    .Q(sig00000441)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056f (
    .C(clk),
    .CE(sig00000002),
    .D(b[50]),
    .Q(sig00000443)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000570 (
    .C(clk),
    .CE(sig00000002),
    .D(b[51]),
    .Q(sig00000444)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000571 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000008b9),
    .Q(sig000003e0)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000572 (
    .I0(sig0000064e),
    .I1(sig0000064f),
    .O(sig00000666)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000573 (
    .I0(sig0000064c),
    .I1(sig0000064d),
    .O(sig00000665)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000574 (
    .I0(b[52]),
    .I1(a[52]),
    .O(sig000008b9)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000575 (
    .I0(b[63]),
    .I1(a[63]),
    .O(sig000005ee)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000576 (
    .I0(a[62]),
    .I1(b[62]),
    .O(sig00000585)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000577 (
    .I0(b[31]),
    .I1(b[30]),
    .I2(a[30]),
    .I3(a[31]),
    .O(sig0000053f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000578 (
    .I0(b[62]),
    .I1(a[62]),
    .O(sig00000595)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000579 (
    .I0(b[62]),
    .I1(a[62]),
    .O(sig00000565)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000057a (
    .I0(b[48]),
    .I1(b[49]),
    .I2(b[50]),
    .I3(b[51]),
    .O(sig00000498)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000057b (
    .I0(a[48]),
    .I1(a[49]),
    .I2(a[50]),
    .I3(a[51]),
    .O(sig00000482)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000057c (
    .I0(b[30]),
    .I1(a[30]),
    .I2(b[31]),
    .I3(a[31]),
    .O(sig0000054f)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000057d (
    .I0(b[61]),
    .I1(b[60]),
    .I2(a[60]),
    .I3(a[61]),
    .O(sig00000584)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000057e (
    .I0(b[29]),
    .I1(b[28]),
    .I2(a[28]),
    .I3(a[29]),
    .O(sig0000053e)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000057f (
    .I0(b[60]),
    .I1(a[60]),
    .I2(b[61]),
    .I3(a[61]),
    .O(sig00000594)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000580 (
    .I0(b[28]),
    .I1(a[28]),
    .I2(b[29]),
    .I3(a[29]),
    .O(sig0000054e)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000581 (
    .I0(b[42]),
    .I1(b[43]),
    .I2(b[44]),
    .I3(b[45]),
    .I4(b[46]),
    .I5(b[47]),
    .O(sig00000497)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000582 (
    .I0(a[42]),
    .I1(a[43]),
    .I2(a[44]),
    .I3(a[45]),
    .I4(a[46]),
    .I5(a[47]),
    .O(sig00000481)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000583 (
    .I0(b[59]),
    .I1(a[59]),
    .I2(b[60]),
    .I3(a[60]),
    .I4(b[61]),
    .I5(a[61]),
    .O(sig0000056e)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000584 (
    .I0(b[59]),
    .I1(b[58]),
    .I2(a[58]),
    .I3(a[59]),
    .O(sig00000583)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000585 (
    .I0(b[27]),
    .I1(b[26]),
    .I2(a[26]),
    .I3(a[27]),
    .O(sig0000053d)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000586 (
    .I0(b[58]),
    .I1(a[58]),
    .I2(b[59]),
    .I3(a[59]),
    .O(sig00000593)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000587 (
    .I0(b[26]),
    .I1(a[26]),
    .I2(b[27]),
    .I3(a[27]),
    .O(sig0000054d)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000588 (
    .I0(b[36]),
    .I1(b[37]),
    .I2(b[38]),
    .I3(b[39]),
    .I4(b[40]),
    .I5(b[41]),
    .O(sig00000496)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000589 (
    .I0(a[36]),
    .I1(a[37]),
    .I2(a[38]),
    .I3(a[39]),
    .I4(a[40]),
    .I5(a[41]),
    .O(sig00000480)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000058a (
    .I0(b[56]),
    .I1(a[56]),
    .I2(b[57]),
    .I3(a[57]),
    .I4(b[58]),
    .I5(a[58]),
    .O(sig0000056d)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000058b (
    .I0(b[57]),
    .I1(b[56]),
    .I2(a[56]),
    .I3(a[57]),
    .O(sig00000582)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000058c (
    .I0(b[25]),
    .I1(b[24]),
    .I2(a[24]),
    .I3(a[25]),
    .O(sig0000053c)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000058d (
    .I0(b[56]),
    .I1(a[56]),
    .I2(b[57]),
    .I3(a[57]),
    .O(sig00000592)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000058e (
    .I0(b[24]),
    .I1(a[24]),
    .I2(b[25]),
    .I3(a[25]),
    .O(sig0000054c)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000058f (
    .I0(b[30]),
    .I1(b[31]),
    .I2(b[32]),
    .I3(b[33]),
    .I4(b[34]),
    .I5(b[35]),
    .O(sig00000495)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000590 (
    .I0(a[30]),
    .I1(a[31]),
    .I2(a[32]),
    .I3(a[33]),
    .I4(a[34]),
    .I5(a[35]),
    .O(sig0000047f)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000591 (
    .I0(b[53]),
    .I1(a[53]),
    .I2(b[54]),
    .I3(a[54]),
    .I4(b[55]),
    .I5(a[55]),
    .O(sig0000056c)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000592 (
    .I0(b[55]),
    .I1(b[54]),
    .I2(a[54]),
    .I3(a[55]),
    .O(sig00000581)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000593 (
    .I0(b[23]),
    .I1(b[22]),
    .I2(a[22]),
    .I3(a[23]),
    .O(sig0000053b)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000594 (
    .I0(sig00000897),
    .I1(sig0000067a),
    .O(sig00000675)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000595 (
    .I0(sig000004cf),
    .I1(sig0000051a),
    .O(sig000005d6)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000596 (
    .I0(sig000004de),
    .I1(sig000004dd),
    .O(sig000005ba)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000597 (
    .I0(sig00000454),
    .I1(sig0000046c),
    .O(sig000005a5)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk00000598 (
    .I0(sig00000486),
    .I1(sig00000470),
    .O(sig000008bc)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk00000599 (
    .I0(sig0000035a),
    .I1(sig0000035d),
    .O(sig000003df)
  );
  LUT2 #(
    .INIT ( 4'h7 ))
  blk0000059a (
    .I0(sig00000320),
    .I1(sig0000001d),
    .O(sig00000143)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000059b (
    .I0(sig0000046c),
    .I1(sig00000454),
    .O(sig000005aa)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk0000059c (
    .I0(sig0000001d),
    .I1(sig00000350),
    .I2(sig0000034f),
    .O(sig00000147)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk0000059d (
    .I0(sig0000001d),
    .I1(sig0000034b),
    .I2(sig0000034a),
    .O(sig00000146)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk0000059e (
    .I0(sig0000001d),
    .I1(sig00000347),
    .I2(sig00000346),
    .O(sig00000145)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk0000059f (
    .I0(sig0000001d),
    .I1(sig00000343),
    .I2(sig00000341),
    .O(sig00000144)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a0 (
    .I0(sig0000001d),
    .I1(sig0000033e),
    .I2(sig0000033d),
    .O(sig00000150)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a1 (
    .I0(sig0000001d),
    .I1(sig0000033a),
    .I2(sig00000339),
    .O(sig0000014f)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a2 (
    .I0(sig0000001d),
    .I1(sig00000335),
    .I2(sig00000334),
    .O(sig0000014e)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a3 (
    .I0(sig0000001d),
    .I1(sig00000331),
    .I2(sig00000330),
    .O(sig0000014d)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a4 (
    .I0(sig0000001d),
    .I1(sig0000032d),
    .I2(sig0000032b),
    .O(sig0000014c)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a5 (
    .I0(sig0000001d),
    .I1(sig00000328),
    .I2(sig00000327),
    .O(sig0000014b)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a6 (
    .I0(sig0000001d),
    .I1(sig00000324),
    .I2(sig00000323),
    .O(sig0000014a)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a7 (
    .I0(sig0000001d),
    .I1(sig00000354),
    .I2(sig00000353),
    .O(sig00000149)
  );
  LUT3 #(
    .INIT ( 8'h57 ))
  blk000005a8 (
    .I0(sig0000001d),
    .I1(sig00000342),
    .I2(sig00000337),
    .O(sig00000148)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000005a9 (
    .I0(sig00000059),
    .I1(sig00000096),
    .I2(sig00000095),
    .O(sig000000c8)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000005aa (
    .I0(sig00000058),
    .I1(sig00000096),
    .I2(sig00000095),
    .O(sig000000c7)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000005ab (
    .I0(sig00000057),
    .I1(sig00000096),
    .I2(sig00000095),
    .O(sig000000c6)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000005ac (
    .I0(sig00000056),
    .I1(sig00000096),
    .I2(sig00000095),
    .O(sig000000c5)
  );
  LUT4 #(
    .INIT ( 16'hA8AA ))
  blk000005ad (
    .I0(sig000004d8),
    .I1(sig000004de),
    .I2(sig000004dd),
    .I3(sig0000046d),
    .O(sig000005eb)
  );
  LUT4 #(
    .INIT ( 16'h22F2 ))
  blk000005ae (
    .I0(sig0000046f),
    .I1(sig000005a6),
    .I2(sig00000485),
    .I3(sig000005ac),
    .O(sig000005a9)
  );
  LUT4 #(
    .INIT ( 16'hF888 ))
  blk000005af (
    .I0(sig00000485),
    .I1(sig000005ac),
    .I2(sig0000046f),
    .I3(sig000005a6),
    .O(sig000005a7)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk000005b0 (
    .I0(sig00000485),
    .I1(sig000005ac),
    .I2(sig0000046f),
    .I3(sig000005a6),
    .O(sig000005a4)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b1 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000351),
    .I3(sig0000033f),
    .O(sig000000ed)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b2 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000350),
    .I3(sig0000033e),
    .O(sig000000ec)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b3 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig0000034f),
    .I3(sig0000033d),
    .O(sig000000eb)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b4 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig0000034e),
    .I3(sig0000033c),
    .O(sig000000ea)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b5 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig0000034c),
    .I3(sig0000033b),
    .O(sig000000e9)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b6 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig0000034b),
    .I3(sig0000033a),
    .O(sig000000e8)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b7 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig0000034a),
    .I3(sig00000339),
    .O(sig000000e7)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b8 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000349),
    .I3(sig00000338),
    .O(sig000000e6)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005b9 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000348),
    .I3(sig00000336),
    .O(sig000000e5)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005ba (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000347),
    .I3(sig00000335),
    .O(sig000000e3)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005bb (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000346),
    .I3(sig00000334),
    .O(sig000000e2)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005bc (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000345),
    .I3(sig00000333),
    .O(sig000000e1)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005bd (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000344),
    .I3(sig00000332),
    .O(sig000000e0)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005be (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000343),
    .I3(sig00000331),
    .O(sig000000df)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005bf (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000341),
    .I3(sig00000330),
    .O(sig000000de)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005c0 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000340),
    .I3(sig0000032f),
    .O(sig000000dd)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005c1 (
    .I0(sig00000096),
    .I1(sig00000095),
    .I2(sig00000059),
    .I3(sig00000055),
    .O(sig000000c4)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005c2 (
    .I0(sig00000096),
    .I1(sig00000095),
    .I2(sig00000058),
    .I3(sig00000053),
    .O(sig000000c2)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005c3 (
    .I0(sig00000096),
    .I1(sig00000095),
    .I2(sig00000057),
    .I3(sig00000052),
    .O(sig000000c1)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk000005c4 (
    .I0(sig00000096),
    .I1(sig00000095),
    .I2(sig00000056),
    .I3(sig00000051),
    .O(sig000000c0)
  );
  LUT4 #(
    .INIT ( 16'hEC4C ))
  blk000005c5 (
    .I0(sig0000046f),
    .I1(sig0000046c),
    .I2(sig000005a6),
    .I3(sig00000454),
    .O(sig000005a8)
  );
  LUT5 #(
    .INIT ( 32'h55555554 ))
  blk000005c6 (
    .I0(sig000004dd),
    .I1(sig0000046d),
    .I2(sig000004de),
    .I3(sig00000528),
    .I4(sig0000051b),
    .O(sig000005b9)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005c7 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000343),
    .I3(sig00000354),
    .I4(sig00000331),
    .O(sig00000104)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005c8 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000341),
    .I3(sig00000353),
    .I4(sig00000330),
    .O(sig00000103)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005c9 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000340),
    .I3(sig00000352),
    .I4(sig0000032f),
    .O(sig00000102)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005ca (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000351),
    .I3(sig0000032e),
    .I4(sig0000033f),
    .O(sig000000dc)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005cb (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000350),
    .I3(sig0000032d),
    .I4(sig0000033e),
    .O(sig000000db)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005cc (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034f),
    .I3(sig0000032b),
    .I4(sig0000033d),
    .O(sig000000da)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005cd (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034e),
    .I3(sig0000032a),
    .I4(sig0000033c),
    .O(sig000000d8)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005ce (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034c),
    .I3(sig00000329),
    .I4(sig0000033b),
    .O(sig000000d7)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005cf (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034b),
    .I3(sig00000328),
    .I4(sig0000033a),
    .O(sig000000d6)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d0 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034a),
    .I3(sig00000327),
    .I4(sig00000339),
    .O(sig000000d5)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d1 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000349),
    .I3(sig00000326),
    .I4(sig00000338),
    .O(sig000000d4)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d2 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000348),
    .I3(sig00000325),
    .I4(sig00000336),
    .O(sig000000d3)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d3 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000347),
    .I3(sig00000324),
    .I4(sig00000335),
    .O(sig000000d2)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d4 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000346),
    .I3(sig00000323),
    .I4(sig00000334),
    .O(sig000000d1)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d5 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000345),
    .I3(sig00000322),
    .I4(sig00000333),
    .O(sig000000d0)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d6 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000344),
    .I3(sig00000355),
    .I4(sig00000332),
    .O(sig000000cf)
  );
  LUT5 #(
    .INIT ( 32'hEC64A820 ))
  blk000005d7 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000339),
    .I3(sig0000034a),
    .I4(sig00000327),
    .O(sig000000ce)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d8 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000059),
    .I3(sig00000050),
    .I4(sig00000055),
    .O(sig000000bf)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005d9 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000058),
    .I3(sig0000004f),
    .I4(sig00000053),
    .O(sig000000be)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005da (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000057),
    .I3(sig0000004e),
    .I4(sig00000052),
    .O(sig000000bd)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk000005db (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000056),
    .I3(sig0000004d),
    .I4(sig00000051),
    .O(sig000000bc)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFF55555554 ))
  blk000005dc (
    .I0(sig000004dd),
    .I1(sig0000046d),
    .I2(sig0000051c),
    .I3(sig00000528),
    .I4(sig0000051b),
    .I5(sig000004de),
    .O(sig000005ed)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAAAAAABAA ))
  blk000005dd (
    .I0(sig000004dd),
    .I1(sig000004de),
    .I2(sig0000046d),
    .I3(sig0000051c),
    .I4(sig00000528),
    .I5(sig0000051b),
    .O(sig000005ec)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk000005de (
    .I0(sig0000046d),
    .I1(sig0000051c),
    .I2(sig00000528),
    .I3(sig0000051b),
    .I4(sig000004dd),
    .I5(sig000004de),
    .O(sig000004ec)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005df (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000351),
    .I3(sig0000033f),
    .I4(sig0000034d),
    .I5(sig0000032e),
    .O(sig00000101)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e0 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig00000350),
    .I3(sig0000033e),
    .I4(sig00000342),
    .I5(sig0000032d),
    .O(sig00000100)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e1 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034f),
    .I3(sig0000033d),
    .I4(sig00000337),
    .I5(sig0000032b),
    .O(sig000000fa)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e2 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034e),
    .I3(sig0000033c),
    .I4(sig0000032c),
    .I5(sig0000032a),
    .O(sig000000ef)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e3 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034c),
    .I3(sig0000033b),
    .I4(sig00000321),
    .I5(sig00000329),
    .O(sig000000e4)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e4 (
    .I0(sig00000021),
    .I1(sig00000022),
    .I2(sig0000034b),
    .I3(sig0000033a),
    .I4(sig00000320),
    .I5(sig00000328),
    .O(sig000000d9)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e5 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000035),
    .I3(sig00000030),
    .I4(sig0000005d),
    .I5(sig0000002c),
    .O(sig000000cd)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e6 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000034),
    .I3(sig0000002f),
    .I4(sig0000005c),
    .I5(sig0000002b),
    .O(sig000000cc)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e7 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000032),
    .I3(sig0000002e),
    .I4(sig0000005b),
    .I5(sig0000002a),
    .O(sig000000cb)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e8 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000031),
    .I3(sig0000002d),
    .I4(sig0000005a),
    .I5(sig00000029),
    .O(sig000000ca)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005e9 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000030),
    .I3(sig0000002c),
    .I4(sig00000054),
    .I5(sig0000005d),
    .O(sig000000c9)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005ea (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000002f),
    .I3(sig0000002b),
    .I4(sig00000049),
    .I5(sig0000005c),
    .O(sig000000c3)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005eb (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000059),
    .I3(sig00000055),
    .I4(sig0000004c),
    .I5(sig00000050),
    .O(sig000000bb)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005ec (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000058),
    .I3(sig00000053),
    .I4(sig0000004b),
    .I5(sig0000004f),
    .O(sig000000ba)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005ed (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000057),
    .I3(sig00000052),
    .I4(sig0000004a),
    .I5(sig0000004e),
    .O(sig000000b9)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005ee (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000002e),
    .I3(sig0000002a),
    .I4(sig0000003e),
    .I5(sig0000005b),
    .O(sig000000b8)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005ef (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000056),
    .I3(sig00000051),
    .I4(sig00000048),
    .I5(sig0000004d),
    .O(sig000000b7)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f0 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000055),
    .I3(sig00000050),
    .I4(sig00000047),
    .I5(sig0000004c),
    .O(sig000000b6)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f1 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000053),
    .I3(sig0000004f),
    .I4(sig00000046),
    .I5(sig0000004b),
    .O(sig000000b5)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f2 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000052),
    .I3(sig0000004e),
    .I4(sig00000045),
    .I5(sig0000004a),
    .O(sig000000b4)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f3 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000051),
    .I3(sig0000004d),
    .I4(sig00000044),
    .I5(sig00000048),
    .O(sig000000b3)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f4 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000050),
    .I3(sig0000004c),
    .I4(sig00000043),
    .I5(sig00000047),
    .O(sig000000b2)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f5 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000004f),
    .I3(sig0000004b),
    .I4(sig00000042),
    .I5(sig00000046),
    .O(sig000000b1)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f6 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000004e),
    .I3(sig0000004a),
    .I4(sig00000041),
    .I5(sig00000045),
    .O(sig000000b0)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f7 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000004d),
    .I3(sig00000048),
    .I4(sig00000040),
    .I5(sig00000044),
    .O(sig000000af)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f8 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000004c),
    .I3(sig00000047),
    .I4(sig0000003f),
    .I5(sig00000043),
    .O(sig000000ae)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005f9 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000002d),
    .I3(sig00000029),
    .I4(sig00000033),
    .I5(sig0000005a),
    .O(sig000000ad)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005fa (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000004b),
    .I3(sig00000046),
    .I4(sig0000003d),
    .I5(sig00000042),
    .O(sig000000ac)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005fb (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000004a),
    .I3(sig00000045),
    .I4(sig0000003c),
    .I5(sig00000041),
    .O(sig000000ab)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005fc (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000048),
    .I3(sig00000044),
    .I4(sig0000003b),
    .I5(sig00000040),
    .O(sig000000aa)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005fd (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000047),
    .I3(sig00000043),
    .I4(sig0000003a),
    .I5(sig0000003f),
    .O(sig000000a9)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005fe (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000046),
    .I3(sig00000042),
    .I4(sig00000039),
    .I5(sig0000003d),
    .O(sig000000a8)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk000005ff (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000045),
    .I3(sig00000041),
    .I4(sig00000038),
    .I5(sig0000003c),
    .O(sig000000a7)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000600 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000044),
    .I3(sig00000040),
    .I4(sig00000037),
    .I5(sig0000003b),
    .O(sig000000a6)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000601 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000043),
    .I3(sig0000003f),
    .I4(sig00000036),
    .I5(sig0000003a),
    .O(sig000000a5)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000602 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000042),
    .I3(sig0000003d),
    .I4(sig00000035),
    .I5(sig00000039),
    .O(sig000000a4)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000603 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000041),
    .I3(sig0000003c),
    .I4(sig00000034),
    .I5(sig00000038),
    .O(sig000000a3)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000604 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000002c),
    .I3(sig0000005d),
    .I4(sig00000028),
    .I5(sig00000054),
    .O(sig000000a2)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000605 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000040),
    .I3(sig0000003b),
    .I4(sig00000032),
    .I5(sig00000037),
    .O(sig000000a1)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000606 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000003f),
    .I3(sig0000003a),
    .I4(sig00000031),
    .I5(sig00000036),
    .O(sig000000a0)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000607 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000003d),
    .I3(sig00000039),
    .I4(sig00000030),
    .I5(sig00000035),
    .O(sig0000009f)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000608 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000003c),
    .I3(sig00000038),
    .I4(sig0000002f),
    .I5(sig00000034),
    .O(sig0000009e)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000609 (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000003b),
    .I3(sig00000037),
    .I4(sig0000002e),
    .I5(sig00000032),
    .O(sig0000009d)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk0000060a (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000003a),
    .I3(sig00000036),
    .I4(sig0000002d),
    .I5(sig00000031),
    .O(sig0000009c)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk0000060b (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000039),
    .I3(sig00000035),
    .I4(sig0000002c),
    .I5(sig00000030),
    .O(sig0000009b)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk0000060c (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000038),
    .I3(sig00000034),
    .I4(sig0000002b),
    .I5(sig0000002f),
    .O(sig0000009a)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk0000060d (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000037),
    .I3(sig00000032),
    .I4(sig0000002a),
    .I5(sig0000002e),
    .O(sig00000099)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk0000060e (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig00000036),
    .I3(sig00000031),
    .I4(sig00000029),
    .I5(sig0000002d),
    .O(sig00000098)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk0000060f (
    .I0(sig00000095),
    .I1(sig00000096),
    .I2(sig0000002b),
    .I3(sig0000005c),
    .I4(sig00000027),
    .I5(sig00000049),
    .O(sig00000097)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000610 (
    .I0(b[54]),
    .I1(a[54]),
    .I2(b[55]),
    .I3(a[55]),
    .O(sig00000591)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000611 (
    .I0(b[22]),
    .I1(a[22]),
    .I2(b[23]),
    .I3(a[23]),
    .O(sig0000054b)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000612 (
    .I0(b[24]),
    .I1(b[25]),
    .I2(b[26]),
    .I3(b[27]),
    .I4(b[28]),
    .I5(b[29]),
    .O(sig00000494)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000613 (
    .I0(a[24]),
    .I1(a[25]),
    .I2(a[26]),
    .I3(a[27]),
    .I4(a[28]),
    .I5(a[29]),
    .O(sig0000047e)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000614 (
    .I0(b[50]),
    .I1(a[50]),
    .I2(b[51]),
    .I3(a[51]),
    .I4(b[52]),
    .I5(a[52]),
    .O(sig0000056b)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000615 (
    .I0(b[53]),
    .I1(b[52]),
    .I2(a[52]),
    .I3(a[53]),
    .O(sig00000580)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000616 (
    .I0(b[21]),
    .I1(b[20]),
    .I2(a[20]),
    .I3(a[21]),
    .O(sig0000053a)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000617 (
    .I0(b[52]),
    .I1(a[52]),
    .I2(b[53]),
    .I3(a[53]),
    .O(sig00000590)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000618 (
    .I0(b[20]),
    .I1(a[20]),
    .I2(b[21]),
    .I3(a[21]),
    .O(sig0000054a)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000619 (
    .I0(b[18]),
    .I1(b[19]),
    .I2(b[20]),
    .I3(b[21]),
    .I4(b[22]),
    .I5(b[23]),
    .O(sig00000493)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000061a (
    .I0(a[18]),
    .I1(a[19]),
    .I2(a[20]),
    .I3(a[21]),
    .I4(a[22]),
    .I5(a[23]),
    .O(sig0000047d)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000061b (
    .I0(b[47]),
    .I1(a[47]),
    .I2(b[48]),
    .I3(a[48]),
    .I4(b[49]),
    .I5(a[49]),
    .O(sig0000056a)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000061c (
    .I0(b[51]),
    .I1(b[50]),
    .I2(a[50]),
    .I3(a[51]),
    .O(sig0000058e)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000061d (
    .I0(b[19]),
    .I1(b[18]),
    .I2(a[18]),
    .I3(a[19]),
    .O(sig00000548)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000061e (
    .I0(b[50]),
    .I1(a[50]),
    .I2(b[51]),
    .I3(a[51]),
    .O(sig0000059e)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000061f (
    .I0(b[18]),
    .I1(a[18]),
    .I2(b[19]),
    .I3(a[19]),
    .O(sig00000558)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000620 (
    .I0(b[12]),
    .I1(b[13]),
    .I2(b[14]),
    .I3(b[15]),
    .I4(b[16]),
    .I5(b[17]),
    .O(sig00000492)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000621 (
    .I0(a[12]),
    .I1(a[13]),
    .I2(a[14]),
    .I3(a[15]),
    .I4(a[16]),
    .I5(a[17]),
    .O(sig0000047c)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000622 (
    .I0(b[44]),
    .I1(a[44]),
    .I2(b[45]),
    .I3(a[45]),
    .I4(b[46]),
    .I5(a[46]),
    .O(sig00000569)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000623 (
    .I0(b[49]),
    .I1(b[48]),
    .I2(a[48]),
    .I3(a[49]),
    .O(sig0000058d)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000624 (
    .I0(b[17]),
    .I1(b[16]),
    .I2(a[16]),
    .I3(a[17]),
    .O(sig00000547)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk00000625 (
    .I0(b[57]),
    .I1(b[56]),
    .I2(b[55]),
    .I3(b[54]),
    .I4(b[53]),
    .I5(b[52]),
    .O(sig00000008)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000626 (
    .I0(b[62]),
    .I1(b[61]),
    .I2(b[60]),
    .I3(b[59]),
    .I4(b[58]),
    .I5(sig00000008),
    .O(sig0000049a)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000627 (
    .I0(b[57]),
    .I1(b[56]),
    .I2(b[55]),
    .I3(b[54]),
    .I4(b[53]),
    .I5(b[52]),
    .O(sig00000013)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000628 (
    .I0(b[62]),
    .I1(b[61]),
    .I2(b[60]),
    .I3(b[59]),
    .I4(b[58]),
    .I5(sig00000013),
    .O(sig00000499)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk00000629 (
    .I0(a[57]),
    .I1(a[56]),
    .I2(a[55]),
    .I3(a[54]),
    .I4(a[53]),
    .I5(a[52]),
    .O(sig0000001a)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000062a (
    .I0(a[62]),
    .I1(a[61]),
    .I2(a[60]),
    .I3(a[59]),
    .I4(a[58]),
    .I5(sig0000001a),
    .O(sig00000484)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk0000062b (
    .I0(a[57]),
    .I1(a[56]),
    .I2(a[55]),
    .I3(a[54]),
    .I4(a[53]),
    .I5(a[52]),
    .O(sig0000001b)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk0000062c (
    .I0(a[62]),
    .I1(a[61]),
    .I2(a[60]),
    .I3(a[59]),
    .I4(a[58]),
    .I5(sig0000001b),
    .O(sig00000483)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000062d (
    .I0(b[48]),
    .I1(a[48]),
    .I2(b[49]),
    .I3(a[49]),
    .O(sig0000059d)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000062e (
    .I0(b[16]),
    .I1(a[16]),
    .I2(b[17]),
    .I3(a[17]),
    .O(sig00000557)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000062f (
    .I0(b[6]),
    .I1(b[7]),
    .I2(b[8]),
    .I3(b[9]),
    .I4(b[10]),
    .I5(b[11]),
    .O(sig00000491)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000630 (
    .I0(a[6]),
    .I1(a[7]),
    .I2(a[8]),
    .I3(a[9]),
    .I4(a[10]),
    .I5(a[11]),
    .O(sig0000047b)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000631 (
    .I0(b[41]),
    .I1(a[41]),
    .I2(b[42]),
    .I3(a[42]),
    .I4(b[43]),
    .I5(a[43]),
    .O(sig00000568)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000632 (
    .I0(b[47]),
    .I1(b[46]),
    .I2(a[46]),
    .I3(a[47]),
    .O(sig0000058c)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000633 (
    .I0(b[15]),
    .I1(b[14]),
    .I2(a[14]),
    .I3(a[15]),
    .O(sig00000546)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000634 (
    .I0(b[46]),
    .I1(a[46]),
    .I2(b[47]),
    .I3(a[47]),
    .O(sig0000059c)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000635 (
    .I0(b[14]),
    .I1(a[14]),
    .I2(b[15]),
    .I3(a[15]),
    .O(sig00000556)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000636 (
    .I0(b[0]),
    .I1(b[1]),
    .I2(b[2]),
    .I3(b[3]),
    .I4(b[4]),
    .I5(b[5]),
    .O(sig00000490)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000637 (
    .I0(a[0]),
    .I1(a[1]),
    .I2(a[2]),
    .I3(a[3]),
    .I4(a[4]),
    .I5(a[5]),
    .O(sig0000047a)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000638 (
    .I0(b[38]),
    .I1(a[38]),
    .I2(b[39]),
    .I3(a[39]),
    .I4(b[40]),
    .I5(a[40]),
    .O(sig00000567)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000639 (
    .I0(b[45]),
    .I1(b[44]),
    .I2(a[44]),
    .I3(a[45]),
    .O(sig0000058b)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000063a (
    .I0(b[13]),
    .I1(b[12]),
    .I2(a[12]),
    .I3(a[13]),
    .O(sig00000545)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000063b (
    .I0(b[44]),
    .I1(a[44]),
    .I2(b[45]),
    .I3(a[45]),
    .O(sig0000059b)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000063c (
    .I0(b[12]),
    .I1(a[12]),
    .I2(b[13]),
    .I3(a[13]),
    .O(sig00000555)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000063d (
    .I0(b[35]),
    .I1(a[35]),
    .I2(b[36]),
    .I3(a[36]),
    .I4(b[37]),
    .I5(a[37]),
    .O(sig00000566)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000063e (
    .I0(b[43]),
    .I1(b[42]),
    .I2(a[42]),
    .I3(a[43]),
    .O(sig0000058a)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000063f (
    .I0(b[11]),
    .I1(b[10]),
    .I2(a[10]),
    .I3(a[11]),
    .O(sig00000544)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000640 (
    .I0(b[42]),
    .I1(a[42]),
    .I2(b[43]),
    .I3(a[43]),
    .O(sig0000059a)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000641 (
    .I0(b[10]),
    .I1(a[10]),
    .I2(b[11]),
    .I3(a[11]),
    .O(sig00000554)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000642 (
    .I0(b[32]),
    .I1(a[32]),
    .I2(b[33]),
    .I3(a[33]),
    .I4(b[34]),
    .I5(a[34]),
    .O(sig00000564)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000643 (
    .I0(sig00000458),
    .I1(sig00000457),
    .O(sig0000035f)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000644 (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e3),
    .O(sig000008a4)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000645 (
    .I0(b[41]),
    .I1(b[40]),
    .I2(a[40]),
    .I3(a[41]),
    .O(sig00000589)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000646 (
    .I0(b[9]),
    .I1(b[8]),
    .I2(a[8]),
    .I3(a[9]),
    .O(sig00000543)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000647 (
    .I0(b[40]),
    .I1(a[40]),
    .I2(b[41]),
    .I3(a[41]),
    .O(sig00000599)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000648 (
    .I0(b[8]),
    .I1(a[8]),
    .I2(b[9]),
    .I3(a[9]),
    .O(sig00000553)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000649 (
    .I0(b[39]),
    .I1(b[38]),
    .I2(a[38]),
    .I3(a[39]),
    .O(sig00000588)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000064a (
    .I0(b[7]),
    .I1(b[6]),
    .I2(a[6]),
    .I3(a[7]),
    .O(sig00000542)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000064b (
    .I0(b[38]),
    .I1(a[38]),
    .I2(b[39]),
    .I3(a[39]),
    .O(sig00000598)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000064c (
    .I0(b[6]),
    .I1(a[6]),
    .I2(b[7]),
    .I3(a[7]),
    .O(sig00000552)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000064d (
    .I0(b[37]),
    .I1(b[36]),
    .I2(a[36]),
    .I3(a[37]),
    .O(sig00000587)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk0000064e (
    .I0(b[5]),
    .I1(b[4]),
    .I2(a[4]),
    .I3(a[5]),
    .O(sig00000541)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000064f (
    .I0(b[36]),
    .I1(a[36]),
    .I2(b[37]),
    .I3(a[37]),
    .O(sig00000597)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000650 (
    .I0(b[4]),
    .I1(a[4]),
    .I2(b[5]),
    .I3(a[5]),
    .O(sig00000551)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000651 (
    .I0(sig0000067d),
    .I1(sig00000897),
    .O(sig00000653)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000652 (
    .I0(sig0000064c),
    .I1(sig0000062f),
    .I2(sig0000062d),
    .O(sig00000660)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000653 (
    .I0(sig0000064c),
    .I1(sig0000062e),
    .I2(sig0000062c),
    .O(sig0000065f)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000654 (
    .I0(sig0000067d),
    .I1(sig00000680),
    .I2(sig0000067c),
    .O(sig00000652)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000655 (
    .I0(sig0000067d),
    .I1(sig0000067f),
    .I2(sig0000067b),
    .O(sig00000651)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000656 (
    .I0(sig0000067d),
    .I1(sig0000067e),
    .I2(sig00000676),
    .O(sig00000650)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000657 (
    .I0(sig00000678),
    .I1(sig00000677),
    .O(sig00000656)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000658 (
    .I0(sig0000064e),
    .I1(sig00000633),
    .I2(sig00000631),
    .O(sig00000662)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000659 (
    .I0(sig0000064e),
    .I1(sig00000632),
    .I2(sig00000630),
    .O(sig00000661)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000065a (
    .I0(sig00000678),
    .I1(sig0000067a),
    .I2(sig00000682),
    .O(sig00000655)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000065b (
    .I0(sig00000678),
    .I1(sig00000679),
    .I2(sig00000681),
    .O(sig00000654)
  );
  LUT5 #(
    .INIT ( 32'h01010100 ))
  blk0000065c (
    .I0(sig00000678),
    .I1(sig000005f1),
    .I2(sig000005f2),
    .I3(sig00000625),
    .I4(sig00000626),
    .O(sig00000643)
  );
  LUT5 #(
    .INIT ( 32'h11110010 ))
  blk0000065d (
    .I0(sig00000678),
    .I1(sig000005f2),
    .I2(sig00000625),
    .I3(sig00000626),
    .I4(sig000005f1),
    .O(sig00000642)
  );
  LUT5 #(
    .INIT ( 32'h01010100 ))
  blk0000065e (
    .I0(sig00000678),
    .I1(sig000005f5),
    .I2(sig000005f6),
    .I3(sig000005f3),
    .I4(sig000005f4),
    .O(sig00000641)
  );
  LUT5 #(
    .INIT ( 32'h11110010 ))
  blk0000065f (
    .I0(sig00000678),
    .I1(sig000005f6),
    .I2(sig000005f3),
    .I3(sig000005f4),
    .I4(sig000005f5),
    .O(sig00000640)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000660 (
    .I0(b[35]),
    .I1(b[34]),
    .I2(a[34]),
    .I3(a[35]),
    .O(sig00000586)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000661 (
    .I0(b[3]),
    .I1(b[2]),
    .I2(a[2]),
    .I3(a[3]),
    .O(sig00000540)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000662 (
    .I0(b[34]),
    .I1(a[34]),
    .I2(b[35]),
    .I3(a[35]),
    .O(sig00000596)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000663 (
    .I0(b[2]),
    .I1(a[2]),
    .I2(b[3]),
    .I3(a[3]),
    .O(sig00000550)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000664 (
    .I0(b[33]),
    .I1(b[32]),
    .I2(a[32]),
    .I3(a[33]),
    .O(sig0000057f)
  );
  LUT4 #(
    .INIT ( 16'h08AE ))
  blk00000665 (
    .I0(b[1]),
    .I1(b[0]),
    .I2(a[0]),
    .I3(a[1]),
    .O(sig00000539)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000666 (
    .I0(b[32]),
    .I1(a[32]),
    .I2(b[33]),
    .I3(a[33]),
    .O(sig0000058f)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000667 (
    .I0(b[0]),
    .I1(a[0]),
    .I2(b[1]),
    .I3(a[1]),
    .O(sig00000549)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk00000668 (
    .I0(sig0000034f),
    .I1(sig00000350),
    .I2(sig00000351),
    .O(sig00000117)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000669 (
    .I0(sig000002a0),
    .I1(sig00000225),
    .I2(sig00000224),
    .I3(sig00000223),
    .O(sig0000068e)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000066a (
    .I0(sig00000226),
    .I1(sig0000021e),
    .I2(sig00000213),
    .I3(sig00000212),
    .O(sig00000687)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000066b (
    .I0(sig000002b7),
    .I1(sig000002b6),
    .I2(sig000002ac),
    .I3(sig000002a1),
    .O(sig0000068d)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000066c (
    .I0(sig0000022a),
    .I1(sig00000229),
    .I2(sig00000228),
    .I3(sig00000227),
    .O(sig00000686)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000066d (
    .I0(sig0000034a),
    .I1(sig0000034b),
    .I2(sig0000034c),
    .I3(sig0000034e),
    .O(sig00000116)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000066e (
    .I0(sig000002bb),
    .I1(sig000002ba),
    .I2(sig000002b9),
    .I3(sig000002b8),
    .O(sig0000068c)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000066f (
    .I0(sig00000215),
    .I1(sig00000214),
    .I2(sig0000022c),
    .I3(sig0000022b),
    .O(sig00000685)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000670 (
    .I0(sig00000346),
    .I1(sig00000347),
    .I2(sig00000348),
    .I3(sig00000349),
    .O(sig00000115)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000671 (
    .I0(sig000002a4),
    .I1(sig000002a3),
    .I2(sig000002a2),
    .I3(sig000002bc),
    .O(sig0000068b)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000672 (
    .I0(sig00000219),
    .I1(sig00000218),
    .I2(sig00000217),
    .I3(sig00000216),
    .O(sig00000684)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000673 (
    .I0(sig00000341),
    .I1(sig00000343),
    .I2(sig00000344),
    .I3(sig00000345),
    .O(sig00000114)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000674 (
    .I0(sig0000021d),
    .I1(sig0000021c),
    .I2(sig0000021b),
    .I3(sig0000021a),
    .O(sig00000690)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000675 (
    .I0(sig000002a8),
    .I1(sig000002a7),
    .I2(sig000002a6),
    .I3(sig000002a5),
    .O(sig0000068a)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000676 (
    .I0(sig0000033d),
    .I1(sig0000033e),
    .I2(sig0000033f),
    .I3(sig00000340),
    .O(sig00000120)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000677 (
    .I0(sig00000222),
    .I1(sig00000221),
    .I2(sig00000220),
    .I3(sig0000021f),
    .O(sig0000068f)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000678 (
    .I0(sig000002ad),
    .I1(sig000002ab),
    .I2(sig000002aa),
    .I3(sig000002a9),
    .O(sig00000689)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000679 (
    .I0(sig00000339),
    .I1(sig0000033a),
    .I2(sig0000033b),
    .I3(sig0000033c),
    .O(sig0000011f)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk0000067a (
    .I0(sig00000603),
    .I1(sig00000601),
    .I2(sig00000600),
    .I3(sig00000602),
    .O(sig00000003)
  );
  LUT6 #(
    .INIT ( 64'h01010100ABABABAA ))
  blk0000067b (
    .I0(sig0000067d),
    .I1(sig00000614),
    .I2(sig00000615),
    .I3(sig00000612),
    .I4(sig00000613),
    .I5(sig00000003),
    .O(sig0000063b)
  );
  LUT4 #(
    .INIT ( 16'hBBAB ))
  blk0000067c (
    .I0(sig00000603),
    .I1(sig00000602),
    .I2(sig00000600),
    .I3(sig00000601),
    .O(sig00000004)
  );
  LUT6 #(
    .INIT ( 64'h05050100AFAFABAA ))
  blk0000067d (
    .I0(sig0000067d),
    .I1(sig00000613),
    .I2(sig00000615),
    .I3(sig00000612),
    .I4(sig00000614),
    .I5(sig00000004),
    .O(sig0000063a)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk0000067e (
    .I0(sig00000608),
    .I1(sig00000605),
    .I2(sig00000604),
    .I3(sig00000607),
    .O(sig00000005)
  );
  LUT6 #(
    .INIT ( 64'h01010100ABABABAA ))
  blk0000067f (
    .I0(sig0000067d),
    .I1(sig00000618),
    .I2(sig00000619),
    .I3(sig00000616),
    .I4(sig00000617),
    .I5(sig00000005),
    .O(sig00000639)
  );
  LUT4 #(
    .INIT ( 16'hBBAB ))
  blk00000680 (
    .I0(sig00000608),
    .I1(sig00000607),
    .I2(sig00000604),
    .I3(sig00000605),
    .O(sig00000006)
  );
  LUT6 #(
    .INIT ( 64'h05050100AFAFABAA ))
  blk00000681 (
    .I0(sig0000067d),
    .I1(sig00000617),
    .I2(sig00000619),
    .I3(sig00000616),
    .I4(sig00000618),
    .I5(sig00000006),
    .O(sig00000638)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk00000682 (
    .I0(sig0000060c),
    .I1(sig0000060a),
    .I2(sig00000609),
    .I3(sig0000060b),
    .O(sig00000007)
  );
  LUT6 #(
    .INIT ( 64'h01010100ABABABAA ))
  blk00000683 (
    .I0(sig0000067d),
    .I1(sig0000061d),
    .I2(sig0000061e),
    .I3(sig0000061a),
    .I4(sig0000061b),
    .I5(sig00000007),
    .O(sig00000637)
  );
  LUT4 #(
    .INIT ( 16'hBBAB ))
  blk00000684 (
    .I0(sig0000060c),
    .I1(sig0000060b),
    .I2(sig00000609),
    .I3(sig0000060a),
    .O(sig00000009)
  );
  LUT6 #(
    .INIT ( 64'h05050100AFAFABAA ))
  blk00000685 (
    .I0(sig0000067d),
    .I1(sig0000061b),
    .I2(sig0000061e),
    .I3(sig0000061a),
    .I4(sig0000061d),
    .I5(sig00000009),
    .O(sig00000636)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk00000686 (
    .I0(sig00000610),
    .I1(sig0000060e),
    .I2(sig0000060d),
    .I3(sig0000060f),
    .O(sig0000000a)
  );
  LUT6 #(
    .INIT ( 64'h01010100ABABABAA ))
  blk00000687 (
    .I0(sig0000067d),
    .I1(sig00000621),
    .I2(sig00000622),
    .I3(sig0000061f),
    .I4(sig00000620),
    .I5(sig0000000a),
    .O(sig00000635)
  );
  LUT4 #(
    .INIT ( 16'hBBAB ))
  blk00000688 (
    .I0(sig00000610),
    .I1(sig0000060f),
    .I2(sig0000060d),
    .I3(sig0000060e),
    .O(sig0000000b)
  );
  LUT6 #(
    .INIT ( 64'h05050100AFAFABAA ))
  blk00000689 (
    .I0(sig0000067d),
    .I1(sig00000620),
    .I2(sig00000622),
    .I3(sig0000061f),
    .I4(sig00000621),
    .I5(sig0000000b),
    .O(sig00000634)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk0000068a (
    .I0(sig000005f9),
    .I1(sig000005f8),
    .I2(sig000005f7),
    .I3(sig000005fa),
    .O(sig0000000c)
  );
  LUT6 #(
    .INIT ( 64'h0202020057575755 ))
  blk0000068b (
    .I0(sig00000678),
    .I1(sig000005fb),
    .I2(sig00000606),
    .I3(sig000005f0),
    .I4(sig000005ef),
    .I5(sig0000000c),
    .O(sig0000063f)
  );
  LUT4 #(
    .INIT ( 16'hBBAB ))
  blk0000068c (
    .I0(sig000005fa),
    .I1(sig000005f9),
    .I2(sig000005f7),
    .I3(sig000005f8),
    .O(sig0000000d)
  );
  LUT6 #(
    .INIT ( 64'h0A0A02005F5F5755 ))
  blk0000068d (
    .I0(sig00000678),
    .I1(sig000005f0),
    .I2(sig00000606),
    .I3(sig000005ef),
    .I4(sig000005fb),
    .I5(sig0000000d),
    .O(sig0000063e)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk0000068e (
    .I0(sig000005fe),
    .I1(sig000005fd),
    .I2(sig000005fc),
    .I3(sig000005ff),
    .O(sig0000000e)
  );
  LUT6 #(
    .INIT ( 64'h0202020057575755 ))
  blk0000068f (
    .I0(sig00000678),
    .I1(sig00000623),
    .I2(sig00000624),
    .I3(sig0000061c),
    .I4(sig00000611),
    .I5(sig0000000e),
    .O(sig0000063d)
  );
  LUT4 #(
    .INIT ( 16'hBBAB ))
  blk00000690 (
    .I0(sig000005ff),
    .I1(sig000005fe),
    .I2(sig000005fc),
    .I3(sig000005fd),
    .O(sig0000000f)
  );
  LUT6 #(
    .INIT ( 64'h0A0A02005F5F5755 ))
  blk00000691 (
    .I0(sig00000678),
    .I1(sig0000061c),
    .I2(sig00000624),
    .I3(sig00000611),
    .I4(sig00000623),
    .I5(sig0000000f),
    .O(sig0000063c)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000692 (
    .I0(sig000002b1),
    .I1(sig000002b0),
    .I2(sig000002af),
    .I3(sig000002ae),
    .O(sig00000688)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000693 (
    .I0(sig00000334),
    .I1(sig00000335),
    .I2(sig00000336),
    .I3(sig00000338),
    .O(sig0000011e)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000694 (
    .I0(sig00000486),
    .I1(sig00000470),
    .O(sig000008bb)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000695 (
    .I0(sig000005a1),
    .I1(sig0000059f),
    .I2(sig000005a0),
    .O(sig000008ba)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000696 (
    .I0(sig0000064e),
    .I1(sig0000064c),
    .I2(sig0000064d),
    .O(sig00000895)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk00000697 (
    .I0(sig000006c7),
    .I1(sig00000695),
    .I2(sig00000699),
    .I3(sig0000069e),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000735)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk00000698 (
    .I0(sig000006c6),
    .I1(sig00000694),
    .I2(sig00000698),
    .I3(sig0000069d),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000734)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk00000699 (
    .I0(sig000006c5),
    .I1(sig00000693),
    .I2(sig00000697),
    .I3(sig0000069b),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000733)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk0000069a (
    .I0(sig000006c4),
    .I1(sig00000692),
    .I2(sig00000696),
    .I3(sig0000069a),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000732)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk0000069b (
    .I0(sig000006bd),
    .I1(sig000006c7),
    .I2(sig00000695),
    .I3(sig00000699),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000731)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk0000069c (
    .I0(sig000006b2),
    .I1(sig000006c6),
    .I2(sig00000694),
    .I3(sig00000698),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000072a)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000069d (
    .I0(sig000006ba),
    .I1(sig000006b6),
    .I2(sig000006bf),
    .I3(sig000006c3),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000723)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000069e (
    .I0(sig000006b9),
    .I1(sig000006b5),
    .I2(sig000006be),
    .I3(sig000006c2),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000722)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000069f (
    .I0(sig000006b8),
    .I1(sig000006b4),
    .I2(sig000006bc),
    .I3(sig000006c1),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000721)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a0 (
    .I0(sig000006b7),
    .I1(sig000006b3),
    .I2(sig000006bb),
    .I3(sig000006c0),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000720)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006a1 (
    .I0(sig000006a7),
    .I1(sig000006c5),
    .I2(sig00000693),
    .I3(sig00000697),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000071f)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a2 (
    .I0(sig000006b6),
    .I1(sig000006b1),
    .I2(sig000006ba),
    .I3(sig000006bf),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000071e)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a3 (
    .I0(sig000006b5),
    .I1(sig000006b0),
    .I2(sig000006b9),
    .I3(sig000006be),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000071d)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a4 (
    .I0(sig000006b4),
    .I1(sig000006af),
    .I2(sig000006b8),
    .I3(sig000006bc),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000071c)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a5 (
    .I0(sig000006b3),
    .I1(sig000006ae),
    .I2(sig000006b7),
    .I3(sig000006bb),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000071b)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a6 (
    .I0(sig000006b1),
    .I1(sig000006ad),
    .I2(sig000006b6),
    .I3(sig000006ba),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000071a)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a7 (
    .I0(sig000006b0),
    .I1(sig000006ac),
    .I2(sig000006b5),
    .I3(sig000006b9),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000719)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a8 (
    .I0(sig000006af),
    .I1(sig000006ab),
    .I2(sig000006b4),
    .I3(sig000006b8),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000718)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006a9 (
    .I0(sig000006ae),
    .I1(sig000006aa),
    .I2(sig000006b3),
    .I3(sig000006b7),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000717)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006aa (
    .I0(sig000006ad),
    .I1(sig000006a9),
    .I2(sig000006b1),
    .I3(sig000006b6),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000716)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ab (
    .I0(sig000006ac),
    .I1(sig000006a8),
    .I2(sig000006b0),
    .I3(sig000006b5),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000715)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006ac (
    .I0(sig0000069c),
    .I1(sig000006c4),
    .I2(sig00000692),
    .I3(sig00000696),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000714)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ad (
    .I0(sig000006ab),
    .I1(sig000006a6),
    .I2(sig000006af),
    .I3(sig000006b4),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000713)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ae (
    .I0(sig000006aa),
    .I1(sig000006a5),
    .I2(sig000006ae),
    .I3(sig000006b3),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000712)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006af (
    .I0(sig000006a9),
    .I1(sig000006a4),
    .I2(sig000006ad),
    .I3(sig000006b1),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000711)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b0 (
    .I0(sig000006a8),
    .I1(sig000006a3),
    .I2(sig000006ac),
    .I3(sig000006b0),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000710)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b1 (
    .I0(sig000006a6),
    .I1(sig000006a2),
    .I2(sig000006ab),
    .I3(sig000006af),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000070f)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b2 (
    .I0(sig000006a5),
    .I1(sig000006a1),
    .I2(sig000006aa),
    .I3(sig000006ae),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000070e)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b3 (
    .I0(sig000006a4),
    .I1(sig000006a0),
    .I2(sig000006a9),
    .I3(sig000006ad),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000070d)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b4 (
    .I0(sig000006a3),
    .I1(sig0000069f),
    .I2(sig000006a8),
    .I3(sig000006ac),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000070c)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b5 (
    .I0(sig000006a2),
    .I1(sig0000069e),
    .I2(sig000006a6),
    .I3(sig000006ab),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000070b)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b6 (
    .I0(sig000006a1),
    .I1(sig0000069d),
    .I2(sig000006a5),
    .I3(sig000006aa),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig0000070a)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006b7 (
    .I0(sig00000691),
    .I1(sig000006bd),
    .I2(sig000006c7),
    .I3(sig00000695),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000709)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b8 (
    .I0(sig000006a0),
    .I1(sig0000069b),
    .I2(sig000006a4),
    .I3(sig000006a9),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000708)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006b9 (
    .I0(sig0000069f),
    .I1(sig0000069a),
    .I2(sig000006a3),
    .I3(sig000006a8),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000707)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ba (
    .I0(sig0000069e),
    .I1(sig00000699),
    .I2(sig000006a2),
    .I3(sig000006a6),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000706)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006bb (
    .I0(sig0000069d),
    .I1(sig00000698),
    .I2(sig000006a1),
    .I3(sig000006a5),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000705)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006bc (
    .I0(sig0000069b),
    .I1(sig00000697),
    .I2(sig000006a0),
    .I3(sig000006a4),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000704)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006bd (
    .I0(sig0000069a),
    .I1(sig00000696),
    .I2(sig0000069f),
    .I3(sig000006a3),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000703)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006be (
    .I0(sig00000699),
    .I1(sig00000695),
    .I2(sig0000069e),
    .I3(sig000006a2),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000702)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006bf (
    .I0(sig00000694),
    .I1(sig00000698),
    .I2(sig0000069d),
    .I3(sig000006a1),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000701)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006c0 (
    .I0(sig00000693),
    .I1(sig00000697),
    .I2(sig0000069b),
    .I3(sig000006a0),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig00000700)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006c1 (
    .I0(sig00000692),
    .I1(sig00000696),
    .I2(sig0000069a),
    .I3(sig0000069f),
    .I4(sig0000064d),
    .I5(sig00000895),
    .O(sig000006ff)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006c2 (
    .I0(sig00000413),
    .I1(sig00000447),
    .I2(sig00000448),
    .I3(sig00000414),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003dc)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006c3 (
    .I0(sig00000412),
    .I1(sig00000446),
    .I2(sig00000447),
    .I3(sig00000413),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003db)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006c4 (
    .I0(sig00000411),
    .I1(sig00000445),
    .I2(sig00000446),
    .I3(sig00000412),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003da)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006c5 (
    .I0(sig0000040e),
    .I1(sig00000442),
    .I2(sig00000445),
    .I3(sig00000411),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d9)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006c6 (
    .I0(sig00000403),
    .I1(sig00000437),
    .I2(sig00000442),
    .I3(sig0000040e),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d8)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006c7 (
    .I0(sig0000040f),
    .I1(sig00000443),
    .I2(sig00000444),
    .I3(sig00000410),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d6)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006c8 (
    .I0(sig0000040d),
    .I1(sig00000441),
    .I2(sig00000443),
    .I3(sig0000040f),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d5)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006c9 (
    .I0(sig000003f8),
    .I1(sig0000042c),
    .I2(sig00000437),
    .I3(sig00000403),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d4)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ca (
    .I0(sig0000040c),
    .I1(sig00000440),
    .I2(sig00000441),
    .I3(sig0000040d),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d3)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006cb (
    .I0(sig0000040b),
    .I1(sig0000043f),
    .I2(sig00000440),
    .I3(sig0000040c),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d2)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006cc (
    .I0(sig0000040a),
    .I1(sig0000043e),
    .I2(sig0000043f),
    .I3(sig0000040b),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d1)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006cd (
    .I0(sig00000409),
    .I1(sig0000043d),
    .I2(sig0000043e),
    .I3(sig0000040a),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003d0)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ce (
    .I0(sig00000408),
    .I1(sig0000043c),
    .I2(sig0000043d),
    .I3(sig00000409),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003cf)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006cf (
    .I0(sig00000407),
    .I1(sig0000043b),
    .I2(sig0000043c),
    .I3(sig00000408),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003ce)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d0 (
    .I0(sig00000406),
    .I1(sig0000043a),
    .I2(sig0000043b),
    .I3(sig00000407),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003cd)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d1 (
    .I0(sig00000405),
    .I1(sig00000439),
    .I2(sig0000043a),
    .I3(sig00000406),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003cc)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d2 (
    .I0(sig00000404),
    .I1(sig00000438),
    .I2(sig00000439),
    .I3(sig00000405),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003cb)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d3 (
    .I0(sig00000402),
    .I1(sig00000436),
    .I2(sig00000438),
    .I3(sig00000404),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003ca)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d4 (
    .I0(sig000003ed),
    .I1(sig00000421),
    .I2(sig0000042c),
    .I3(sig000003f8),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c9)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d5 (
    .I0(sig00000401),
    .I1(sig00000435),
    .I2(sig00000436),
    .I3(sig00000402),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c8)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d6 (
    .I0(sig00000400),
    .I1(sig00000434),
    .I2(sig00000435),
    .I3(sig00000401),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c7)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d7 (
    .I0(sig000003ff),
    .I1(sig00000433),
    .I2(sig00000434),
    .I3(sig00000400),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c6)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d8 (
    .I0(sig000003fe),
    .I1(sig00000432),
    .I2(sig00000433),
    .I3(sig000003ff),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c5)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006d9 (
    .I0(sig000003fd),
    .I1(sig00000431),
    .I2(sig00000432),
    .I3(sig000003fe),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c4)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006da (
    .I0(sig000003fc),
    .I1(sig00000430),
    .I2(sig00000431),
    .I3(sig000003fd),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c3)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006db (
    .I0(sig000003fb),
    .I1(sig0000042f),
    .I2(sig00000430),
    .I3(sig000003fc),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c2)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006dc (
    .I0(sig000003fa),
    .I1(sig0000042e),
    .I2(sig0000042f),
    .I3(sig000003fb),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c1)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006dd (
    .I0(sig000003f9),
    .I1(sig0000042d),
    .I2(sig0000042e),
    .I3(sig000003fa),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003c0)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006de (
    .I0(sig000003f7),
    .I1(sig0000042b),
    .I2(sig0000042d),
    .I3(sig000003f9),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003bf)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006df (
    .I0(sig000003e2),
    .I1(sig00000416),
    .I2(sig00000421),
    .I3(sig000003ed),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003be)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e0 (
    .I0(sig000003f6),
    .I1(sig0000042a),
    .I2(sig0000042b),
    .I3(sig000003f7),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003bd)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e1 (
    .I0(sig000003f5),
    .I1(sig00000429),
    .I2(sig0000042a),
    .I3(sig000003f6),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003bc)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e2 (
    .I0(sig000003f4),
    .I1(sig00000428),
    .I2(sig00000429),
    .I3(sig000003f5),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003bb)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e3 (
    .I0(sig000003f3),
    .I1(sig00000427),
    .I2(sig00000428),
    .I3(sig000003f4),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003ba)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e4 (
    .I0(sig000003f2),
    .I1(sig00000426),
    .I2(sig00000427),
    .I3(sig000003f3),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b9)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e5 (
    .I0(sig000003f1),
    .I1(sig00000425),
    .I2(sig00000426),
    .I3(sig000003f2),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b8)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e6 (
    .I0(sig000003f0),
    .I1(sig00000424),
    .I2(sig00000425),
    .I3(sig000003f1),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b7)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e7 (
    .I0(sig000003ef),
    .I1(sig00000423),
    .I2(sig00000424),
    .I3(sig000003f0),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b6)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e8 (
    .I0(sig000003ee),
    .I1(sig00000422),
    .I2(sig00000423),
    .I3(sig000003ef),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b5)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006e9 (
    .I0(sig000003ec),
    .I1(sig00000420),
    .I2(sig00000422),
    .I3(sig000003ee),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b4)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ea (
    .I0(sig000003e1),
    .I1(sig00000415),
    .I2(sig00000416),
    .I3(sig000003e2),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b3)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006eb (
    .I0(sig000003eb),
    .I1(sig0000041f),
    .I2(sig00000420),
    .I3(sig000003ec),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b2)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ec (
    .I0(sig000003ea),
    .I1(sig0000041e),
    .I2(sig0000041f),
    .I3(sig000003eb),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b1)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ed (
    .I0(sig000003e9),
    .I1(sig0000041d),
    .I2(sig0000041e),
    .I3(sig000003ea),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003b0)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ee (
    .I0(sig000003e8),
    .I1(sig0000041c),
    .I2(sig0000041d),
    .I3(sig000003e9),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003af)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006ef (
    .I0(sig000003e7),
    .I1(sig0000041b),
    .I2(sig0000041c),
    .I3(sig000003e8),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003ae)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006f0 (
    .I0(sig000003e6),
    .I1(sig0000041a),
    .I2(sig0000041b),
    .I3(sig000003e7),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003ad)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006f1 (
    .I0(sig000003e5),
    .I1(sig00000419),
    .I2(sig0000041a),
    .I3(sig000003e6),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003ac)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006f2 (
    .I0(sig000003e4),
    .I1(sig00000418),
    .I2(sig00000419),
    .I3(sig000003e5),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003ab)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006f3 (
    .I0(sig000003e3),
    .I1(sig00000417),
    .I2(sig00000418),
    .I3(sig000003e4),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003aa)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk000006f4 (
    .I0(sig00000414),
    .I1(sig00000448),
    .I2(sig00000417),
    .I3(sig000003e3),
    .I4(sig000003e0),
    .I5(sig000008ba),
    .O(sig000003a9)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006f5 (
    .I0(sig0000061a),
    .I1(sig00000609),
    .I2(sig000005f7),
    .I3(sig000005ef),
    .I4(sig00000897),
    .I5(sig00000896),
    .O(sig0000076a)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006f6 (
    .I0(sig0000061b),
    .I1(sig0000060a),
    .I2(sig000005f8),
    .I3(sig000005f0),
    .I4(sig00000897),
    .I5(sig00000896),
    .O(sig00000769)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006f7 (
    .I0(sig0000061d),
    .I1(sig0000060b),
    .I2(sig000005f9),
    .I3(sig000005fb),
    .I4(sig00000897),
    .I5(sig00000896),
    .O(sig00000768)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006f8 (
    .I0(sig0000061e),
    .I1(sig0000060c),
    .I2(sig000005fa),
    .I3(sig00000606),
    .I4(sig00000897),
    .I5(sig00000896),
    .O(sig00000761)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006f9 (
    .I0(sig0000061f),
    .I1(sig0000060d),
    .I2(sig000005fc),
    .I3(sig00000611),
    .I4(sig00000897),
    .I5(sig00000896),
    .O(sig00000756)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006fa (
    .I0(sig00000620),
    .I1(sig0000060e),
    .I2(sig000005fd),
    .I3(sig0000061c),
    .I4(sig00000897),
    .I5(sig00000896),
    .O(sig0000074b)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000006fb (
    .I0(sig00000621),
    .I1(sig0000060f),
    .I2(sig000005fe),
    .I3(sig00000623),
    .I4(sig00000897),
    .I5(sig00000896),
    .O(sig00000740)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000006fc (
    .I0(sig00000021),
    .I1(sig00000022),
    .O(sig000003de)
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  blk000006fd (
    .I0(sig000004b2),
    .I1(sig000004b3),
    .I2(sig000004b0),
    .O(sig000005dd)
  );
  LUT5 #(
    .INIT ( 32'h00008000 ))
  blk000006fe (
    .I0(sig000004b4),
    .I1(sig000004b5),
    .I2(sig000004b6),
    .I3(sig000004ad),
    .I4(sig000004ae),
    .O(sig000005dc)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000006ff (
    .I0(sig000004ac),
    .I1(sig000004af),
    .I2(sig000004b1),
    .I3(sig000004ab),
    .I4(sig000005dd),
    .I5(sig000005dc),
    .O(sig000005db)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000700 (
    .I0(sig000002b5),
    .I1(sig000002b4),
    .I2(sig000002b3),
    .I3(sig000002b2),
    .O(sig00000683)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000701 (
    .I0(sig00000330),
    .I1(sig00000331),
    .I2(sig00000332),
    .I3(sig00000333),
    .O(sig0000011d)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000702 (
    .I0(sig0000032b),
    .I1(sig0000032d),
    .I2(sig0000032e),
    .I3(sig0000032f),
    .O(sig0000011c)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000703 (
    .I0(sig00000327),
    .I1(sig00000328),
    .I2(sig00000329),
    .I3(sig0000032a),
    .O(sig0000011b)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000704 (
    .I0(sig00000323),
    .I1(sig00000324),
    .I2(sig00000325),
    .I3(sig00000326),
    .O(sig0000011a)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000705 (
    .I0(sig00000353),
    .I1(sig00000354),
    .I2(sig00000355),
    .I3(sig00000322),
    .O(sig00000119)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000706 (
    .I0(sig00000337),
    .I1(sig00000342),
    .I2(sig0000034d),
    .I3(sig00000352),
    .O(sig00000118)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk00000707 (
    .I0(sig00000320),
    .I1(sig00000321),
    .I2(sig0000032c),
    .O(sig00000113)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000708 (
    .I0(sig00000458),
    .I1(sig00000460),
    .O(sig00000368)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000709 (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004eb),
    .O(sig000008ad)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000070a (
    .I0(sig00000458),
    .I1(sig0000044b),
    .I2(sig00000463),
    .O(sig000005cc)
  );
  LUT5 #(
    .INIT ( 32'h04FBFB04 ))
  blk0000070b (
    .I0(sig00000156),
    .I1(sig0000020a),
    .I2(sig000002bd),
    .I3(sig000001a3),
    .I4(sig0000029f),
    .O(sig0000030c)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk0000070c (
    .I0(sig0000065e),
    .I1(sig0000065d),
    .I2(sig000006df),
    .I3(sig000006dc),
    .I4(sig000006db),
    .I5(sig000006dd),
    .O(sig0000086f)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk0000070d (
    .I0(sig000001d5),
    .I1(sig00000357),
    .I2(sig00000359),
    .I3(sig00000071),
    .I4(sig0000035e),
    .I5(sig00000073),
    .O(sig000002f1)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000070e (
    .I0(sig00000458),
    .I1(sig0000045f),
    .O(sig00000367)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk0000070f (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004ea),
    .O(sig000008ac)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000710 (
    .I0(sig00000458),
    .I1(sig00000453),
    .I2(sig0000046b),
    .O(sig000005d5)
  );
  LUT5 #(
    .INIT ( 32'h04FBFB04 ))
  blk00000711 (
    .I0(sig00000156),
    .I1(sig00000209),
    .I2(sig000002bd),
    .I3(sig000001a2),
    .I4(sig0000029f),
    .O(sig0000030b)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000712 (
    .I0(sig00000852),
    .I1(sig00000851),
    .I2(sig00000846),
    .I3(sig00000848),
    .I4(sig00000849),
    .I5(sig00000847),
    .O(sig00000889)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000713 (
    .I0(sig0000065e),
    .I1(sig0000065d),
    .I2(sig000006e0),
    .I3(sig000006dd),
    .I4(sig000006dc),
    .I5(sig000006df),
    .O(sig0000086e)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk00000714 (
    .I0(sig000001d4),
    .I1(sig00000357),
    .I2(sig00000359),
    .I3(sig00000070),
    .I4(sig0000035e),
    .I5(sig00000072),
    .O(sig000002f0)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000715 (
    .I0(sig00000458),
    .I1(sig0000045e),
    .O(sig00000366)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000716 (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e9),
    .O(sig000008ab)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000717 (
    .I0(sig00000458),
    .I1(sig00000452),
    .I2(sig0000046a),
    .O(sig000005d4)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000718 (
    .I0(sig00000852),
    .I1(sig00000851),
    .I2(sig00000845),
    .I3(sig00000847),
    .I4(sig00000848),
    .I5(sig00000846),
    .O(sig00000888)
  );
  LUT6 #(
    .INIT ( 64'hF7B3E6A2D591C480 ))
  blk00000719 (
    .I0(sig0000065e),
    .I1(sig0000065d),
    .I2(sig000006e1),
    .I3(sig000006df),
    .I4(sig000006dd),
    .I5(sig000006e0),
    .O(sig0000086d)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk0000071a (
    .I0(sig000001a1),
    .I1(sig0000029f),
    .I2(sig00000156),
    .I3(sig00000208),
    .I4(sig000002bd),
    .I5(sig0000020a),
    .O(sig0000030a)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk0000071b (
    .I0(sig000001d3),
    .I1(sig00000357),
    .I2(sig00000359),
    .I3(sig0000006f),
    .I4(sig0000035e),
    .I5(sig00000071),
    .O(sig000002ef)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000071c (
    .I0(sig00000458),
    .I1(sig0000045d),
    .O(sig00000365)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk0000071d (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e8),
    .O(sig000008aa)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000071e (
    .I0(sig00000458),
    .I1(sig00000451),
    .I2(sig00000469),
    .O(sig000005d3)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk0000071f (
    .I0(sig00000847),
    .I1(sig00000845),
    .I2(sig00000846),
    .I3(sig00000844),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000887)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000720 (
    .I0(sig000006e1),
    .I1(sig000006df),
    .I2(sig000006e0),
    .I3(sig000006e2),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig0000086c)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk00000721 (
    .I0(sig000001a0),
    .I1(sig0000029f),
    .I2(sig00000156),
    .I3(sig00000207),
    .I4(sig000002bd),
    .I5(sig00000209),
    .O(sig00000309)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk00000722 (
    .I0(sig000001d2),
    .I1(sig00000357),
    .I2(sig00000359),
    .I3(sig0000006e),
    .I4(sig0000035e),
    .I5(sig00000070),
    .O(sig000002ee)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000723 (
    .I0(sig00000458),
    .I1(sig0000045c),
    .O(sig00000364)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000724 (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e7),
    .O(sig000008a9)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000725 (
    .I0(sig00000458),
    .I1(sig00000450),
    .I2(sig00000468),
    .O(sig000005d2)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000726 (
    .I0(sig00000844),
    .I1(sig00000846),
    .I2(sig00000845),
    .I3(sig00000843),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000886)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000727 (
    .I0(sig000006e2),
    .I1(sig000006e0),
    .I2(sig000006e1),
    .I3(sig000006e3),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig0000086b)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk00000728 (
    .I0(sig0000019f),
    .I1(sig0000029f),
    .I2(sig00000156),
    .I3(sig00000206),
    .I4(sig000002bd),
    .I5(sig00000208),
    .O(sig00000308)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk00000729 (
    .I0(sig000001d1),
    .I1(sig00000357),
    .I2(sig00000359),
    .I3(sig0000006d),
    .I4(sig0000035e),
    .I5(sig0000006f),
    .O(sig000002ed)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000072a (
    .I0(sig00000458),
    .I1(sig0000045b),
    .O(sig00000363)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk0000072b (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e6),
    .O(sig000008a8)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000072c (
    .I0(sig00000458),
    .I1(sig0000044f),
    .I2(sig00000467),
    .O(sig000005d1)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000072d (
    .I0(sig00000843),
    .I1(sig00000845),
    .I2(sig00000844),
    .I3(sig00000842),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000885)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000072e (
    .I0(sig000006e3),
    .I1(sig000006e1),
    .I2(sig000006e2),
    .I3(sig000006e4),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig0000086a)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk0000072f (
    .I0(sig0000019e),
    .I1(sig0000029f),
    .I2(sig00000156),
    .I3(sig00000205),
    .I4(sig000002bd),
    .I5(sig00000207),
    .O(sig00000307)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk00000730 (
    .I0(sig000001cf),
    .I1(sig00000357),
    .I2(sig00000359),
    .I3(sig0000006c),
    .I4(sig0000035e),
    .I5(sig0000006e),
    .O(sig000002ec)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000731 (
    .I0(sig00000458),
    .I1(sig0000045a),
    .O(sig00000362)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000732 (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e5),
    .O(sig000008a7)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000733 (
    .I0(sig00000458),
    .I1(sig0000044e),
    .I2(sig00000466),
    .O(sig000005d0)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000734 (
    .I0(sig00000842),
    .I1(sig00000844),
    .I2(sig00000843),
    .I3(sig00000841),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000884)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000735 (
    .I0(sig000006e4),
    .I1(sig000006e2),
    .I2(sig000006e3),
    .I3(sig000006e5),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000868)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk00000736 (
    .I0(sig0000019d),
    .I1(sig0000029f),
    .I2(sig00000156),
    .I3(sig00000204),
    .I4(sig000002bd),
    .I5(sig00000206),
    .O(sig00000306)
  );
  LUT6 #(
    .INIT ( 64'h6666999666666966 ))
  blk00000737 (
    .I0(sig000001ce),
    .I1(sig00000357),
    .I2(sig00000359),
    .I3(sig0000006b),
    .I4(sig0000035e),
    .I5(sig0000006d),
    .O(sig000002eb)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000738 (
    .I0(sig00000458),
    .I1(sig00000459),
    .O(sig00000361)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000739 (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e4),
    .O(sig000008a6)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000073a (
    .I0(sig00000458),
    .I1(sig0000044d),
    .I2(sig00000465),
    .O(sig000005cf)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000073b (
    .I0(sig00000841),
    .I1(sig00000843),
    .I2(sig00000842),
    .I3(sig0000083f),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000882)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000073c (
    .I0(sig000006e5),
    .I1(sig000006e3),
    .I2(sig000006e4),
    .I3(sig000006e6),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000867)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000073d (
    .I0(sig0000019c),
    .I1(sig00000205),
    .I2(sig00000203),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000305)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000073e (
    .I0(sig000001cd),
    .I1(sig0000006c),
    .I2(sig00000069),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002ea)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000073f (
    .I0(sig00000458),
    .I1(sig00000456),
    .O(sig00000360)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000740 (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e2),
    .O(sig000008a5)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000741 (
    .I0(sig00000458),
    .I1(sig0000044c),
    .I2(sig00000464),
    .O(sig000005ce)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000742 (
    .I0(sig0000083f),
    .I1(sig00000842),
    .I2(sig00000841),
    .I3(sig0000083e),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000881)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000743 (
    .I0(sig000006e6),
    .I1(sig000006e4),
    .I2(sig000006e5),
    .I3(sig000006e7),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000866)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000744 (
    .I0(sig0000019a),
    .I1(sig00000204),
    .I2(sig00000201),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000303)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000745 (
    .I0(sig000001cc),
    .I1(sig0000006b),
    .I2(sig00000068),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e9)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000746 (
    .I0(sig00000458),
    .I1(sig0000044a),
    .I2(sig00000462),
    .O(sig000005cd)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000747 (
    .I0(sig0000083e),
    .I1(sig00000841),
    .I2(sig0000083f),
    .I3(sig0000083d),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000880)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000748 (
    .I0(sig000006e7),
    .I1(sig000006e5),
    .I2(sig000006e6),
    .I3(sig000006e8),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000865)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000749 (
    .I0(sig00000199),
    .I1(sig00000203),
    .I2(sig00000200),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000302)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000074a (
    .I0(sig000001cb),
    .I1(sig00000069),
    .I2(sig00000067),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e8)
  );
  LUT3 #(
    .INIT ( 8'h20 ))
  blk0000074b (
    .I0(sig0000012e),
    .I1(sig00000095),
    .I2(sig00000141),
    .O(sig00000010)
  );
  LUT5 #(
    .INIT ( 32'h8F808080 ))
  blk0000074c (
    .I0(sig00000124),
    .I1(sig00000136),
    .I2(sig00000095),
    .I3(sig00000123),
    .I4(sig00000135),
    .O(sig00000011)
  );
  LUT3 #(
    .INIT ( 8'hF8 ))
  blk0000074d (
    .I0(sig0000012e),
    .I1(sig00000141),
    .I2(sig00000095),
    .O(sig00000012)
  );
  LUT6 #(
    .INIT ( 64'hFFF8F7F00F080700 ))
  blk0000074e (
    .I0(sig0000012f),
    .I1(sig00000142),
    .I2(sig00000096),
    .I3(sig00000010),
    .I4(sig00000012),
    .I5(sig00000011),
    .O(sig00000153)
  );
  LUT5 #(
    .INIT ( 32'h8F808080 ))
  blk0000074f (
    .I0(sig00000126),
    .I1(sig00000138),
    .I2(sig00000095),
    .I3(sig00000125),
    .I4(sig00000137),
    .O(sig00000014)
  );
  LUT5 #(
    .INIT ( 32'h1DDD3FFF ))
  blk00000750 (
    .I0(sig0000013d),
    .I1(sig00000095),
    .I2(sig0000013e),
    .I3(sig0000012b),
    .I4(sig0000012a),
    .O(sig00000015)
  );
  LUT3 #(
    .INIT ( 8'hDF ))
  blk00000751 (
    .I0(sig0000013f),
    .I1(sig00000095),
    .I2(sig0000012c),
    .O(sig00000016)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000752 (
    .I0(sig00000095),
    .I1(sig0000013f),
    .I2(sig0000012c),
    .O(sig00000017)
  );
  LUT6 #(
    .INIT ( 64'h80F000708FFF0F7F ))
  blk00000753 (
    .I0(sig0000012d),
    .I1(sig00000140),
    .I2(sig00000096),
    .I3(sig00000016),
    .I4(sig00000017),
    .I5(sig00000015),
    .O(sig00000152)
  );
  LUT3 #(
    .INIT ( 8'h1B ))
  blk00000754 (
    .I0(sig00000458),
    .I1(sig00000461),
    .I2(sig00000449),
    .O(sig000005ab)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000755 (
    .I0(sig0000083d),
    .I1(sig0000083f),
    .I2(sig0000083e),
    .I3(sig0000083c),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000087f)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000756 (
    .I0(sig000006e8),
    .I1(sig000006e6),
    .I2(sig000006e7),
    .I3(sig000006ea),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000864)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000757 (
    .I0(sig00000198),
    .I1(sig00000201),
    .I2(sig000001ff),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000301)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000758 (
    .I0(sig000001ca),
    .I1(sig00000068),
    .I2(sig00000066),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e7)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000759 (
    .I0(sig0000083c),
    .I1(sig0000083e),
    .I2(sig0000083d),
    .I3(sig0000083b),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000087e)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000075a (
    .I0(sig000006ea),
    .I1(sig000006e7),
    .I2(sig000006e8),
    .I3(sig000006eb),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000863)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000075b (
    .I0(sig00000197),
    .I1(sig00000200),
    .I2(sig000001fe),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000300)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000075c (
    .I0(sig000001c9),
    .I1(sig00000067),
    .I2(sig00000065),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e6)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000075d (
    .I0(sig0000083b),
    .I1(sig0000083d),
    .I2(sig0000083c),
    .I3(sig0000083a),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000087d)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000075e (
    .I0(sig000006eb),
    .I1(sig000006e8),
    .I2(sig000006ea),
    .I3(sig000006ec),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000862)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000075f (
    .I0(sig00000196),
    .I1(sig000001ff),
    .I2(sig000001fd),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig000002ff)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000760 (
    .I0(sig000001c8),
    .I1(sig00000066),
    .I2(sig00000064),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e5)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000761 (
    .I0(sig0000083a),
    .I1(sig0000083c),
    .I2(sig0000083b),
    .I3(sig00000839),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000087c)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000762 (
    .I0(sig000006ec),
    .I1(sig000006ea),
    .I2(sig000006eb),
    .I3(sig000006ed),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000861)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000763 (
    .I0(sig00000195),
    .I1(sig000001fe),
    .I2(sig000001fc),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig000002fe)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000764 (
    .I0(sig000001c7),
    .I1(sig00000065),
    .I2(sig00000063),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e4)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000765 (
    .I0(sig00000839),
    .I1(sig0000083b),
    .I2(sig0000083a),
    .I3(sig00000838),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000087b)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000766 (
    .I0(sig000006ed),
    .I1(sig000006eb),
    .I2(sig000006ec),
    .I3(sig000006ee),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000860)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000767 (
    .I0(sig00000194),
    .I1(sig000001fd),
    .I2(sig000001fb),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig000002fd)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000768 (
    .I0(sig000001c6),
    .I1(sig00000064),
    .I2(sig00000062),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e3)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000769 (
    .I0(sig00000897),
    .I1(sig00000678),
    .I2(sig0000067d),
    .O(sig00000896)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000076a (
    .I0(sig000004c6),
    .I1(sig0000065b),
    .I2(sig000004c7),
    .I3(sig0000062b),
    .O(sig000005d9)
  );
  LUT5 #(
    .INIT ( 32'h00000009 ))
  blk0000076b (
    .I0(sig000004c8),
    .I1(sig0000062a),
    .I2(sig000004ca),
    .I3(sig000004cb),
    .I4(sig000004c9),
    .O(sig000005da)
  );
  LUT6 #(
    .INIT ( 64'h0000000000009009 ))
  blk0000076c (
    .I0(sig000004c2),
    .I1(sig0000065d),
    .I2(sig000004c3),
    .I3(sig0000065e),
    .I4(sig000004c4),
    .I5(sig000004cc),
    .O(sig000005d8)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000076d (
    .I0(sig00000838),
    .I1(sig0000083a),
    .I2(sig00000839),
    .I3(sig00000837),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000087a)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000076e (
    .I0(sig000006ed),
    .I1(sig000006ec),
    .I2(sig000006ee),
    .I3(sig000006ef),
    .I4(sig0000065e),
    .I5(sig0000065d),
    .O(sig0000085f)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000076f (
    .I0(sig00000193),
    .I1(sig000001fc),
    .I2(sig000001fa),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig000002fc)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000770 (
    .I0(sig000001dc),
    .I1(sig00000063),
    .I2(sig00000061),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e2)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000771 (
    .I0(sig00000837),
    .I1(sig00000839),
    .I2(sig00000838),
    .I3(sig00000836),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000879)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000772 (
    .I0(sig000006ef),
    .I1(sig000006ed),
    .I2(sig000006ee),
    .I3(sig000006f0),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000877)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000773 (
    .I0(sig00000192),
    .I1(sig000001fb),
    .I2(sig000001f9),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig000002fb)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000774 (
    .I0(sig000001db),
    .I1(sig00000062),
    .I2(sig00000060),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e1)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000775 (
    .I0(sig00000837),
    .I1(sig00000838),
    .I2(sig00000836),
    .I3(sig00000850),
    .I4(sig00000852),
    .I5(sig00000851),
    .O(sig00000891)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000776 (
    .I0(sig000006f0),
    .I1(sig000006ee),
    .I2(sig000006ef),
    .I3(sig000006f1),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000876)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000777 (
    .I0(sig00000191),
    .I1(sig000001fa),
    .I2(sig000001f8),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig000002fa)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000778 (
    .I0(sig000001da),
    .I1(sig00000061),
    .I2(sig00000094),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002e0)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000779 (
    .I0(sig00000850),
    .I1(sig00000837),
    .I2(sig00000836),
    .I3(sig0000084f),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000890)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000077a (
    .I0(sig000006f1),
    .I1(sig000006ef),
    .I2(sig000006f0),
    .I3(sig000006f2),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000875)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000077b (
    .I0(sig000001aa),
    .I1(sig000001f9),
    .I2(sig00000211),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000314)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000077c (
    .I0(sig000001d9),
    .I1(sig00000060),
    .I2(sig00000093),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002f8)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000077d (
    .I0(sig0000084f),
    .I1(sig00000836),
    .I2(sig00000850),
    .I3(sig0000084e),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000088f)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000077e (
    .I0(sig000006f2),
    .I1(sig000006f0),
    .I2(sig000006f1),
    .I3(sig000006f3),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000874)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000077f (
    .I0(sig000001a9),
    .I1(sig000001f8),
    .I2(sig00000210),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000313)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000780 (
    .I0(sig000001d8),
    .I1(sig00000094),
    .I2(sig00000092),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002f7)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000781 (
    .I0(sig0000084e),
    .I1(sig00000850),
    .I2(sig0000084f),
    .I3(sig0000084d),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000088e)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000782 (
    .I0(sig000006f3),
    .I1(sig000006f1),
    .I2(sig000006f2),
    .I3(sig000006f5),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000873)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000783 (
    .I0(sig000001a8),
    .I1(sig00000211),
    .I2(sig0000020f),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000312)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000784 (
    .I0(sig000001d7),
    .I1(sig00000093),
    .I2(sig00000091),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002f6)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000785 (
    .I0(sig0000084d),
    .I1(sig0000084f),
    .I2(sig0000084e),
    .I3(sig0000084c),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000088d)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk00000786 (
    .I0(sig000006f5),
    .I1(sig000006f2),
    .I2(sig000006f3),
    .I3(sig000006f6),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000872)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000787 (
    .I0(sig000001a7),
    .I1(sig00000210),
    .I2(sig0000020e),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000311)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000788 (
    .I0(sig000001d6),
    .I1(sig00000092),
    .I2(sig0000008b),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002f5)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000789 (
    .I0(sig0000049c),
    .I1(sig0000049b),
    .I2(sig000004e1),
    .O(sig000008a3)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000078a (
    .I0(sig0000084c),
    .I1(sig0000084e),
    .I2(sig0000084d),
    .I3(sig0000084b),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000088c)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000078b (
    .I0(sig000006f6),
    .I1(sig000006f3),
    .I2(sig000006f5),
    .I3(sig000006f7),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000871)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000078c (
    .I0(sig000001a6),
    .I1(sig0000020f),
    .I2(sig0000020d),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000310)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk0000078d (
    .I0(sig000001d0),
    .I1(sig00000091),
    .I2(sig00000080),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002f4)
  );
  LUT6 #(
    .INIT ( 64'hFF00AAAAF0F0CCCC ))
  blk0000078e (
    .I0(sig0000084b),
    .I1(sig0000084d),
    .I2(sig0000084c),
    .I3(sig0000084a),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000088b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000078f (
    .I0(sig000006f5),
    .I1(sig000006f6),
    .I2(sig000006f7),
    .I3(sig000006f8),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000870)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000790 (
    .I0(sig000001a5),
    .I1(sig0000020e),
    .I2(sig0000020c),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig0000030f)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000791 (
    .I0(sig000001c5),
    .I1(sig0000008b),
    .I2(sig00000075),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002f3)
  );
  LUT6 #(
    .INIT ( 64'hAAAACCCCFF00F0F0 ))
  blk00000792 (
    .I0(sig00000840),
    .I1(sig0000084a),
    .I2(sig0000084c),
    .I3(sig0000084b),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig0000088a)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk00000793 (
    .I0(sig000006f6),
    .I1(sig000006f8),
    .I2(sig000006f7),
    .I3(sig000006f9),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000869)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000794 (
    .I0(sig000001a4),
    .I1(sig0000020d),
    .I2(sig0000020b),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig0000030e)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000795 (
    .I0(sig000001c4),
    .I1(sig00000080),
    .I2(sig0000006a),
    .I3(sig0000035e),
    .I4(sig00000359),
    .I5(sig00000357),
    .O(sig000002f2)
  );
  LUT5 #(
    .INIT ( 32'hF30CF50A ))
  blk00000796 (
    .I0(sig0000005f),
    .I1(sig00000075),
    .I2(sig0000035e),
    .I3(sig00000357),
    .I4(sig00000359),
    .O(sig000002c2)
  );
  LUT6 #(
    .INIT ( 64'hAAAACCCCFF00F0F0 ))
  blk00000797 (
    .I0(sig00000835),
    .I1(sig00000840),
    .I2(sig0000084b),
    .I3(sig0000084a),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000883)
  );
  LUT6 #(
    .INIT ( 64'hAAAACCCCFF00F0F0 ))
  blk00000798 (
    .I0(sig000006fa),
    .I1(sig000006f9),
    .I2(sig000006f7),
    .I3(sig000006f8),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig0000085e)
  );
  LUT6 #(
    .INIT ( 64'h559955A5AA66AA5A ))
  blk00000799 (
    .I0(sig0000019b),
    .I1(sig0000020c),
    .I2(sig00000202),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig0000030d)
  );
  LUT5 #(
    .INIT ( 32'hF30CF50A ))
  blk0000079a (
    .I0(sig0000005e),
    .I1(sig0000006a),
    .I2(sig0000035e),
    .I3(sig00000357),
    .I4(sig00000359),
    .O(sig000002c1)
  );
  LUT6 #(
    .INIT ( 64'hAAAACCCCF0F0FF00 ))
  blk0000079b (
    .I0(sig00000834),
    .I1(sig00000835),
    .I2(sig00000840),
    .I3(sig0000084a),
    .I4(sig00000851),
    .I5(sig00000852),
    .O(sig00000878)
  );
  LUT6 #(
    .INIT ( 64'h33C33399CC3CCC66 ))
  blk0000079c (
    .I0(sig000001f7),
    .I1(sig00000190),
    .I2(sig0000020b),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig00000304)
  );
  LUT6 #(
    .INIT ( 64'h33C33399CC3CCC66 ))
  blk0000079d (
    .I0(sig000001f6),
    .I1(sig0000018f),
    .I2(sig00000202),
    .I3(sig000002bd),
    .I4(sig00000156),
    .I5(sig0000029f),
    .O(sig000002f9)
  );
  LUT5 #(
    .INIT ( 32'h00CCAAF0 ))
  blk0000079e (
    .I0(sig000006fa),
    .I1(sig000006f9),
    .I2(sig000006f8),
    .I3(sig0000065e),
    .I4(sig0000065d),
    .O(sig0000085b)
  );
  LUT4 #(
    .INIT ( 16'hFF51 ))
  blk0000079f (
    .I0(sig000006fa),
    .I1(sig000006f9),
    .I2(sig0000065d),
    .I3(sig0000065e),
    .O(sig0000085a)
  );
  LUT6 #(
    .INIT ( 64'hAAAACCCCFF00F0F0 ))
  blk000007a0 (
    .I0(sig000006fa),
    .I1(sig000006f9),
    .I2(sig000006f7),
    .I3(sig000006f8),
    .I4(sig0000065d),
    .I5(sig0000065e),
    .O(sig00000859)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007a1 (
    .C(clk),
    .D(sig00000002),
    .R(sig000003e0),
    .Q(sig00000351)
  );
  FDS #(
    .INIT ( 1'b0 ))
  blk000007a2 (
    .C(clk),
    .D(sig000003d7),
    .S(sig000003e0),
    .Q(sig00000350)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007a3 (
    .C(clk),
    .D(sig00000385),
    .R(sig000008bb),
    .Q(sig00000173)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007a4 (
    .C(clk),
    .D(sig00000386),
    .R(sig000008bb),
    .Q(sig00000174)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007a5 (
    .C(clk),
    .D(sig00000387),
    .R(sig000008bb),
    .Q(sig0000017f)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007a6 (
    .C(clk),
    .D(sig00000388),
    .R(sig000008bb),
    .Q(sig00000188)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007a7 (
    .C(clk),
    .D(sig00000389),
    .R(sig000008bb),
    .Q(sig00000189)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007a8 (
    .C(clk),
    .D(sig0000038b),
    .R(sig000008bb),
    .Q(sig0000018a)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007a9 (
    .C(clk),
    .D(sig0000038c),
    .R(sig000008bb),
    .Q(sig0000018b)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007aa (
    .C(clk),
    .D(sig0000038d),
    .R(sig000008bb),
    .Q(sig0000018c)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007ab (
    .C(clk),
    .D(sig0000038e),
    .R(sig000008bb),
    .Q(sig0000018d)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007ac (
    .C(clk),
    .D(sig0000038f),
    .R(sig000008bb),
    .Q(sig0000018e)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007ad (
    .C(clk),
    .D(sig00000390),
    .R(sig000008bb),
    .Q(sig00000175)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007ae (
    .C(clk),
    .D(sig00000391),
    .R(sig000008bb),
    .Q(sig00000176)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007af (
    .C(clk),
    .D(sig00000392),
    .R(sig000008bb),
    .Q(sig00000177)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b0 (
    .C(clk),
    .D(sig00000393),
    .R(sig000008bb),
    .Q(sig00000178)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b1 (
    .C(clk),
    .D(sig00000394),
    .R(sig000008bb),
    .Q(sig00000179)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b2 (
    .C(clk),
    .D(sig00000396),
    .R(sig000008bb),
    .Q(sig0000017a)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b3 (
    .C(clk),
    .D(sig00000397),
    .R(sig000008bb),
    .Q(sig0000017b)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b4 (
    .C(clk),
    .D(sig00000398),
    .R(sig000008bb),
    .Q(sig0000017c)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b5 (
    .C(clk),
    .D(sig00000399),
    .R(sig000008bb),
    .Q(sig0000017d)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b6 (
    .C(clk),
    .D(sig0000039a),
    .R(sig000008bb),
    .Q(sig0000017e)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b7 (
    .C(clk),
    .D(sig0000039b),
    .R(sig000008bb),
    .Q(sig00000180)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b8 (
    .C(clk),
    .D(sig0000039c),
    .R(sig000008bb),
    .Q(sig00000181)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007b9 (
    .C(clk),
    .D(sig0000039d),
    .R(sig000008bb),
    .Q(sig00000182)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007ba (
    .C(clk),
    .D(sig0000039e),
    .R(sig000008bb),
    .Q(sig00000183)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007bb (
    .C(clk),
    .D(sig0000039f),
    .R(sig000008bb),
    .Q(sig00000184)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007bc (
    .C(clk),
    .D(sig000003a1),
    .R(sig000008bb),
    .Q(sig00000185)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007bd (
    .C(clk),
    .D(sig000003a2),
    .R(sig000008bb),
    .Q(sig00000186)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007be (
    .C(clk),
    .D(sig00000002),
    .R(sig000008bb),
    .Q(sig00000187)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007bf (
    .C(clk),
    .D(sig00000374),
    .R(sig000008bb),
    .Q(sig000001dd)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c0 (
    .C(clk),
    .D(sig0000037f),
    .R(sig000008bb),
    .Q(sig000001de)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c1 (
    .C(clk),
    .D(sig0000038a),
    .R(sig000008bb),
    .Q(sig000001e9)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c2 (
    .C(clk),
    .D(sig00000395),
    .R(sig000008bb),
    .Q(sig000001ef)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c3 (
    .C(clk),
    .D(sig000003a0),
    .R(sig000008bb),
    .Q(sig000001f0)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c4 (
    .C(clk),
    .D(sig000003a3),
    .R(sig000008bb),
    .Q(sig000001f1)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c5 (
    .C(clk),
    .D(sig000003a4),
    .R(sig000008bb),
    .Q(sig000001f2)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c6 (
    .C(clk),
    .D(sig000003a5),
    .R(sig000008bb),
    .Q(sig000001f3)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c7 (
    .C(clk),
    .D(sig000003a6),
    .R(sig000008bb),
    .Q(sig000001f4)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c8 (
    .C(clk),
    .D(sig000003a7),
    .R(sig000008bb),
    .Q(sig000001f5)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007c9 (
    .C(clk),
    .D(sig00000375),
    .R(sig000008bb),
    .Q(sig000001df)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007ca (
    .C(clk),
    .D(sig00000376),
    .R(sig000008bb),
    .Q(sig000001e0)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007cb (
    .C(clk),
    .D(sig00000377),
    .R(sig000008bb),
    .Q(sig000001e1)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007cc (
    .C(clk),
    .D(sig00000378),
    .R(sig000008bb),
    .Q(sig000001e2)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007cd (
    .C(clk),
    .D(sig00000379),
    .R(sig000008bb),
    .Q(sig000001e3)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007ce (
    .C(clk),
    .D(sig0000037a),
    .R(sig000008bb),
    .Q(sig000001e4)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007cf (
    .C(clk),
    .D(sig0000037b),
    .R(sig000008bb),
    .Q(sig000001e5)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007d0 (
    .C(clk),
    .D(sig0000037c),
    .R(sig000008bb),
    .Q(sig000001e6)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007d1 (
    .C(clk),
    .D(sig0000037d),
    .R(sig000008bb),
    .Q(sig000001e7)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007d2 (
    .C(clk),
    .D(sig0000037e),
    .R(sig000008bb),
    .Q(sig000001e8)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007d3 (
    .C(clk),
    .D(sig00000380),
    .R(sig000008bb),
    .Q(sig000001ea)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007d4 (
    .C(clk),
    .D(sig00000381),
    .R(sig000008bb),
    .Q(sig000001eb)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007d5 (
    .C(clk),
    .D(sig00000382),
    .R(sig000008bb),
    .Q(sig000001ec)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007d6 (
    .C(clk),
    .D(sig00000383),
    .R(sig000008bb),
    .Q(sig000001ed)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk000007d7 (
    .C(clk),
    .D(sig00000384),
    .R(sig000008bb),
    .Q(sig000001ee)
  );
  FDS #(
    .INIT ( 1'b0 ))
  blk000007d8 (
    .C(clk),
    .D(sig000005bf),
    .S(sig000004d1),
    .Q(sig000004e0)
  );
  LUT4 #(
    .INIT ( 16'h1054 ))
  blk000007d9 (
    .I0(sig000004d4),
    .I1(sig000004d0),
    .I2(sig000004d2),
    .I3(sig000004d6),
    .O(sig000005bf)
  );
  FDRS #(
    .INIT ( 1'b0 ))
  blk000007da (
    .C(clk),
    .D(sig000005be),
    .R(sig000004d1),
    .S(sig000004d0),
    .Q(sig000004df)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000007db (
    .I0(sig000004d2),
    .I1(sig000004d4),
    .O(sig000005be)
  );
  LUT5 #(
    .INIT ( 32'hCF8FC080 ))
  blk000007dc (
    .I0(sig00000139),
    .I1(sig00000127),
    .I2(sig00000096),
    .I3(sig00000095),
    .I4(sig00000014),
    .O(sig00000154)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000007dd (
    .I0(sig000002c0),
    .O(sig00000281)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000007de (
    .I0(sig00000130),
    .O(sig0000027f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000007df (
    .I0(sig000004c5),
    .I1(sig0000065c),
    .O(sig00000511)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000007e0 (
    .I0(sig00000894),
    .O(sig00000853)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000007e1 (
    .I0(sig0000085d),
    .O(sig000007fb)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000007e2 (
    .I0(sig0000029f),
    .O(sig00000280)
  );
  LUT4 #(
    .INIT ( 16'h0F09 ))
  blk000007e3 (
    .I0(sig000007f3),
    .I1(sig000004e1),
    .I2(sig0000049c),
    .I3(sig0000049b),
    .O(sig000008a2)
  );
  LUT5 #(
    .INIT ( 32'h8F808080 ))
  blk000007e4 (
    .I0(sig0000013c),
    .I1(sig00000129),
    .I2(sig00000096),
    .I3(sig0000013a),
    .I4(sig00000122),
    .O(sig00000018)
  );
  LUT6 #(
    .INIT ( 64'hFEAEAEAE54040404 ))
  blk000007e5 (
    .I0(sig00000095),
    .I1(sig00000121),
    .I2(sig00000096),
    .I3(sig00000128),
    .I4(sig0000013b),
    .I5(sig00000018),
    .O(sig00000151)
  );
  LUT5 #(
    .INIT ( 32'hFFFFFFFE ))
  blk000007e6 (
    .I0(sig0000001e),
    .I1(sig00000023),
    .I2(sig00000024),
    .I3(sig00000025),
    .I4(sig00000026),
    .O(sig00000019)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFF8F00000 ))
  blk000007e7 (
    .I0(sig0000001c),
    .I1(sig0000001f),
    .I2(sig00000020),
    .I3(sig0000001d),
    .I4(sig000003de),
    .I5(sig00000019),
    .O(sig000003dd)
  );
  LUT5 #(
    .INIT ( 32'h90000000 ))
  blk000007e8 (
    .I0(sig000004c5),
    .I1(sig0000065c),
    .I2(sig000005d9),
    .I3(sig000005da),
    .I4(sig000005d8),
    .O(sig000005d7)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007e9 (
    .I0(sig000006c3),
    .I1(sig0000064d),
    .I2(sig0000064c),
    .O(sig00000730)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007ea (
    .I0(sig000006c2),
    .I1(sig0000064d),
    .I2(sig0000064c),
    .O(sig0000072f)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007eb (
    .I0(sig000006c1),
    .I1(sig0000064d),
    .I2(sig0000064c),
    .O(sig0000072e)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007ec (
    .I0(sig000006c0),
    .I1(sig0000064d),
    .I2(sig0000064c),
    .O(sig0000072d)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007ed (
    .I0(sig000005ef),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000767)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007ee (
    .I0(sig000005f0),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000766)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007ef (
    .I0(sig000005fb),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000765)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f0 (
    .I0(sig00000606),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000764)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f1 (
    .I0(sig00000611),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000763)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f2 (
    .I0(sig0000061c),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000762)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f3 (
    .I0(sig00000623),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000760)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f4 (
    .I0(sig00000624),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig0000075f)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f5 (
    .I0(sig00000625),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig0000075e)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f6 (
    .I0(sig00000626),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig0000075d)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f7 (
    .I0(sig000005f1),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig0000075c)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f8 (
    .I0(sig000005f2),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig0000075b)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007f9 (
    .I0(sig000005f3),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig0000075a)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007fa (
    .I0(sig000005f4),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000759)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007fb (
    .I0(sig000005f5),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000758)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007fc (
    .I0(sig000005f6),
    .I1(sig00000897),
    .I2(sig0000067d),
    .O(sig00000757)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007fd (
    .I0(sig00000351),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000ff)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007fe (
    .I0(sig00000350),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000fe)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk000007ff (
    .I0(sig0000034f),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000fd)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000800 (
    .I0(sig0000034e),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000fc)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000801 (
    .I0(sig0000034c),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000fb)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000802 (
    .I0(sig0000034b),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f9)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000803 (
    .I0(sig0000034a),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f8)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000804 (
    .I0(sig00000349),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f7)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000805 (
    .I0(sig00000348),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f6)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000806 (
    .I0(sig00000347),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f5)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000807 (
    .I0(sig00000346),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f4)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000808 (
    .I0(sig00000345),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f3)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000809 (
    .I0(sig00000344),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f2)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk0000080a (
    .I0(sig00000343),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f1)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk0000080b (
    .I0(sig00000341),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000f0)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk0000080c (
    .I0(sig00000340),
    .I1(sig00000022),
    .I2(sig00000021),
    .O(sig000000ee)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000080d (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005ef),
    .I3(sig000005f7),
    .O(sig00000755)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000080e (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005f0),
    .I3(sig000005f8),
    .O(sig00000754)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000080f (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005fb),
    .I3(sig000005f9),
    .O(sig00000753)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000810 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000606),
    .I3(sig000005fa),
    .O(sig00000752)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000811 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000611),
    .I3(sig000005fc),
    .O(sig00000751)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000812 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig0000061c),
    .I3(sig000005fd),
    .O(sig00000750)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000813 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000623),
    .I3(sig000005fe),
    .O(sig0000074f)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000814 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000624),
    .I3(sig000005ff),
    .O(sig0000074e)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000815 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000625),
    .I3(sig00000600),
    .O(sig0000074d)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000816 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000626),
    .I3(sig00000601),
    .O(sig0000074c)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000817 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005f1),
    .I3(sig00000602),
    .O(sig0000074a)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000818 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005f2),
    .I3(sig00000603),
    .O(sig00000749)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000819 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005f3),
    .I3(sig00000604),
    .O(sig00000748)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000081a (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005f4),
    .I3(sig00000605),
    .O(sig00000747)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000081b (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005f5),
    .I3(sig00000607),
    .O(sig00000746)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000081c (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig000005f6),
    .I3(sig00000608),
    .O(sig00000745)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000081d (
    .I0(sig0000064d),
    .I1(sig0000064c),
    .I2(sig000006c3),
    .I3(sig000006bf),
    .O(sig0000072c)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000081e (
    .I0(sig0000064d),
    .I1(sig0000064c),
    .I2(sig000006c2),
    .I3(sig000006be),
    .O(sig0000072b)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk0000081f (
    .I0(sig0000064d),
    .I1(sig0000064c),
    .I2(sig000006c1),
    .I3(sig000006bc),
    .O(sig00000729)
  );
  LUT4 #(
    .INIT ( 16'h5140 ))
  blk00000820 (
    .I0(sig0000064d),
    .I1(sig0000064c),
    .I2(sig000006c0),
    .I3(sig000006bb),
    .O(sig00000728)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000821 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000046c),
    .I3(sig000005a1),
    .I4(sig00000454),
    .O(sig000005ea)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000822 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000410),
    .I3(sig000005a1),
    .I4(sig00000444),
    .O(sig000003d7)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000823 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000427),
    .I3(sig000005a1),
    .I4(sig000003f3),
    .O(sig00000385)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000824 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000428),
    .I3(sig000005a1),
    .I4(sig000003f4),
    .O(sig00000386)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000825 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000429),
    .I3(sig000005a1),
    .I4(sig000003f5),
    .O(sig00000387)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000826 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000042a),
    .I3(sig000005a1),
    .I4(sig000003f6),
    .O(sig00000388)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000827 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000042b),
    .I3(sig000005a1),
    .I4(sig000003f7),
    .O(sig00000389)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000828 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000042d),
    .I3(sig000005a1),
    .I4(sig000003f9),
    .O(sig0000038b)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000829 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000042e),
    .I3(sig000005a1),
    .I4(sig000003fa),
    .O(sig0000038c)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000082a (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000042f),
    .I3(sig000005a1),
    .I4(sig000003fb),
    .O(sig0000038d)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000082b (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000430),
    .I3(sig000005a1),
    .I4(sig000003fc),
    .O(sig0000038e)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000082c (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000431),
    .I3(sig000005a1),
    .I4(sig000003fd),
    .O(sig0000038f)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000082d (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000432),
    .I3(sig000005a1),
    .I4(sig000003fe),
    .O(sig00000390)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000082e (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000433),
    .I3(sig000005a1),
    .I4(sig000003ff),
    .O(sig00000391)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000082f (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000434),
    .I3(sig000005a1),
    .I4(sig00000400),
    .O(sig00000392)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000830 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000435),
    .I3(sig000005a1),
    .I4(sig00000401),
    .O(sig00000393)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000831 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000436),
    .I3(sig000005a1),
    .I4(sig00000402),
    .O(sig00000394)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000832 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000438),
    .I3(sig000005a1),
    .I4(sig00000404),
    .O(sig00000396)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000833 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000439),
    .I3(sig000005a1),
    .I4(sig00000405),
    .O(sig00000397)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000834 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000043a),
    .I3(sig000005a1),
    .I4(sig00000406),
    .O(sig00000398)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000835 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000043b),
    .I3(sig000005a1),
    .I4(sig00000407),
    .O(sig00000399)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000836 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000043c),
    .I3(sig000005a1),
    .I4(sig00000408),
    .O(sig0000039a)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000837 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000043d),
    .I3(sig000005a1),
    .I4(sig00000409),
    .O(sig0000039b)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000838 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000043e),
    .I3(sig000005a1),
    .I4(sig0000040a),
    .O(sig0000039c)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000839 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000043f),
    .I3(sig000005a1),
    .I4(sig0000040b),
    .O(sig0000039d)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000083a (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000440),
    .I3(sig000005a1),
    .I4(sig0000040c),
    .O(sig0000039e)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000083b (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000441),
    .I3(sig000005a1),
    .I4(sig0000040d),
    .O(sig0000039f)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000083c (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000443),
    .I3(sig000005a1),
    .I4(sig0000040f),
    .O(sig000003a1)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000083d (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000444),
    .I3(sig000005a1),
    .I4(sig00000410),
    .O(sig000003a2)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000083e (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000415),
    .I3(sig000005a1),
    .I4(sig000003e1),
    .O(sig00000374)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000083f (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000416),
    .I3(sig000005a1),
    .I4(sig000003e2),
    .O(sig0000037f)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000840 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000421),
    .I3(sig000005a1),
    .I4(sig000003ed),
    .O(sig0000038a)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000841 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000042c),
    .I3(sig000005a1),
    .I4(sig000003f8),
    .O(sig00000395)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000842 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000437),
    .I3(sig000005a1),
    .I4(sig00000403),
    .O(sig000003a0)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000843 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000442),
    .I3(sig000005a1),
    .I4(sig0000040e),
    .O(sig000003a3)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000844 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000445),
    .I3(sig000005a1),
    .I4(sig00000411),
    .O(sig000003a4)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000845 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000446),
    .I3(sig000005a1),
    .I4(sig00000412),
    .O(sig000003a5)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000846 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000447),
    .I3(sig000005a1),
    .I4(sig00000413),
    .O(sig000003a6)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000847 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000448),
    .I3(sig000005a1),
    .I4(sig00000414),
    .O(sig000003a7)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000848 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000417),
    .I3(sig000005a1),
    .I4(sig000003e3),
    .O(sig00000375)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000849 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000418),
    .I3(sig000005a1),
    .I4(sig000003e4),
    .O(sig00000376)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000084a (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000419),
    .I3(sig000005a1),
    .I4(sig000003e5),
    .O(sig00000377)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000084b (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000041a),
    .I3(sig000005a1),
    .I4(sig000003e6),
    .O(sig00000378)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000084c (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000041b),
    .I3(sig000005a1),
    .I4(sig000003e7),
    .O(sig00000379)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000084d (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000041c),
    .I3(sig000005a1),
    .I4(sig000003e8),
    .O(sig0000037a)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000084e (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000041d),
    .I3(sig000005a1),
    .I4(sig000003e9),
    .O(sig0000037b)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk0000084f (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000041e),
    .I3(sig000005a1),
    .I4(sig000003ea),
    .O(sig0000037c)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000850 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig0000041f),
    .I3(sig000005a1),
    .I4(sig000003eb),
    .O(sig0000037d)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000851 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000420),
    .I3(sig000005a1),
    .I4(sig000003ec),
    .O(sig0000037e)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000852 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000422),
    .I3(sig000005a1),
    .I4(sig000003ee),
    .O(sig00000380)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000853 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000423),
    .I3(sig000005a1),
    .I4(sig000003ef),
    .O(sig00000381)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000854 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000424),
    .I3(sig000005a1),
    .I4(sig000003f0),
    .O(sig00000382)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000855 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000425),
    .I3(sig000005a1),
    .I4(sig000003f1),
    .O(sig00000383)
  );
  LUT5 #(
    .INIT ( 32'hF0F7F080 ))
  blk00000856 (
    .I0(sig000005a0),
    .I1(sig0000059f),
    .I2(sig00000426),
    .I3(sig000005a1),
    .I4(sig000003f2),
    .O(sig00000384)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000857 (
    .I0(sig0000064d),
    .I1(sig0000064c),
    .I2(sig000006ba),
    .I3(sig000006bf),
    .I4(sig0000064e),
    .I5(sig000006c3),
    .O(sig00000727)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000858 (
    .I0(sig0000064d),
    .I1(sig0000064c),
    .I2(sig000006b9),
    .I3(sig000006be),
    .I4(sig0000064e),
    .I5(sig000006c2),
    .O(sig00000726)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000859 (
    .I0(sig0000064d),
    .I1(sig0000064c),
    .I2(sig000006b8),
    .I3(sig000006bc),
    .I4(sig0000064e),
    .I5(sig000006c1),
    .O(sig00000725)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000085a (
    .I0(sig0000064d),
    .I1(sig0000064c),
    .I2(sig000006b7),
    .I3(sig000006bb),
    .I4(sig0000064e),
    .I5(sig000006c0),
    .O(sig00000724)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000085b (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000618),
    .I3(sig00000607),
    .I4(sig00000678),
    .I5(sig000005f5),
    .O(sig0000076c)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000085c (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000619),
    .I3(sig00000608),
    .I4(sig00000678),
    .I5(sig000005f6),
    .O(sig0000076b)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000085d (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000609),
    .I3(sig000005f7),
    .I4(sig00000678),
    .I5(sig000005ef),
    .O(sig00000744)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000085e (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig0000060a),
    .I3(sig000005f8),
    .I4(sig00000678),
    .I5(sig000005f0),
    .O(sig00000743)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000085f (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig0000060b),
    .I3(sig000005f9),
    .I4(sig00000678),
    .I5(sig000005fb),
    .O(sig00000742)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000860 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig0000060c),
    .I3(sig000005fa),
    .I4(sig00000678),
    .I5(sig00000606),
    .O(sig00000741)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000861 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig0000060d),
    .I3(sig000005fc),
    .I4(sig00000678),
    .I5(sig00000611),
    .O(sig0000073f)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000862 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig0000060e),
    .I3(sig000005fd),
    .I4(sig00000678),
    .I5(sig0000061c),
    .O(sig0000073e)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000863 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig0000060f),
    .I3(sig000005fe),
    .I4(sig00000678),
    .I5(sig00000623),
    .O(sig0000073d)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000864 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000610),
    .I3(sig000005ff),
    .I4(sig00000678),
    .I5(sig00000624),
    .O(sig0000073c)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000865 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000612),
    .I3(sig00000600),
    .I4(sig00000678),
    .I5(sig00000625),
    .O(sig0000073b)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000866 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000613),
    .I3(sig00000601),
    .I4(sig00000678),
    .I5(sig00000626),
    .O(sig0000073a)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000867 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000614),
    .I3(sig00000602),
    .I4(sig00000678),
    .I5(sig000005f1),
    .O(sig00000739)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000868 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000615),
    .I3(sig00000603),
    .I4(sig00000678),
    .I5(sig000005f2),
    .O(sig00000738)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000869 (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000616),
    .I3(sig00000604),
    .I4(sig00000678),
    .I5(sig000005f3),
    .O(sig00000737)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000086a (
    .I0(sig00000897),
    .I1(sig0000067d),
    .I2(sig00000617),
    .I3(sig00000605),
    .I4(sig00000678),
    .I5(sig000005f4),
    .O(sig00000736)
  );
  LUT6 #(
    .INIT ( 64'hAAA80200AA882200 ))
  blk0000086b (
    .I0(sig000003e0),
    .I1(sig000005a1),
    .I2(sig0000059f),
    .I3(sig00000415),
    .I4(sig000003e1),
    .I5(sig000005a0),
    .O(sig000003a8)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000086c (
    .I0(sig00000455),
    .O(sig00000316)
  );
  INV   blk0000086d (
    .I(sig000004c4),
    .O(sig0000050f)
  );
  INV   blk0000086e (
    .I(sig000004c9),
    .O(sig00000515)
  );
  INV   blk0000086f (
    .I(sig000004ca),
    .O(sig00000516)
  );
  INV   blk00000870 (
    .I(sig000004cb),
    .O(sig00000517)
  );
  INV   blk00000871 (
    .I(sig000004cc),
    .O(sig00000518)
  );
  LUT6 #(
    .INIT ( 64'hF5F5F4F501010001 ))
  blk00000872 (
    .I0(sig000004d4),
    .I1(sig000004d0),
    .I2(sig000004d1),
    .I3(sig000004d2),
    .I4(sig000004d3),
    .I5(sig000004d5),
    .O(sig000005bc)
  );
  LUT6 #(
    .INIT ( 64'hF5F4F4F401000000 ))
  blk00000873 (
    .I0(sig000004d4),
    .I1(sig000004d0),
    .I2(sig000004d1),
    .I3(sig000004d2),
    .I4(sig000004d3),
    .I5(sig000004d5),
    .O(sig000005bd)
  );
  MUXF7   blk00000874 (
    .I0(sig000005bd),
    .I1(sig000005bc),
    .S(sig000004da),
    .O(sig000005bb)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000875 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000173),
    .Q(sig00000157),
    .Q15(NLW_blk00000875_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000876 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000157),
    .Q(sig0000018f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000877 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000001d),
    .Q(sig00000358),
    .Q15(NLW_blk00000877_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000878 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000358),
    .Q(sig00000359)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000879 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000005a3),
    .Q(sig00000356),
    .Q15(NLW_blk00000879_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000087a (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000356),
    .Q(sig00000357)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000087b (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000174),
    .Q(sig00000158),
    .Q15(NLW_blk0000087b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000087c (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000158),
    .Q(sig00000190)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000087d (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000017f),
    .Q(sig00000163),
    .Q15(NLW_blk0000087d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000087e (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000163),
    .Q(sig0000019b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000087f (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000018a),
    .Q(sig0000016e),
    .Q15(NLW_blk0000087f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000880 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000016e),
    .Q(sig000001a6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000881 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000188),
    .Q(sig0000016c),
    .Q15(NLW_blk00000881_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000882 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000016c),
    .Q(sig000001a4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000883 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000189),
    .Q(sig0000016d),
    .Q15(NLW_blk00000883_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000884 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000016d),
    .Q(sig000001a5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000885 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000018b),
    .Q(sig0000016f),
    .Q15(NLW_blk00000885_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000886 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000016f),
    .Q(sig000001a7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000887 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000018c),
    .Q(sig00000170),
    .Q15(NLW_blk00000887_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000888 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000170),
    .Q(sig000001a8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000889 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000175),
    .Q(sig00000159),
    .Q15(NLW_blk00000889_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000088a (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000159),
    .Q(sig00000191)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000088b (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000018d),
    .Q(sig00000171),
    .Q15(NLW_blk0000088b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000088c (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000171),
    .Q(sig000001a9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000088d (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000018e),
    .Q(sig00000172),
    .Q15(NLW_blk0000088d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000088e (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000172),
    .Q(sig000001aa)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000088f (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000176),
    .Q(sig0000015a),
    .Q15(NLW_blk0000088f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000890 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000015a),
    .Q(sig00000192)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000891 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000177),
    .Q(sig0000015b),
    .Q15(NLW_blk00000891_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000892 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000015b),
    .Q(sig00000193)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000893 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000178),
    .Q(sig0000015c),
    .Q15(NLW_blk00000893_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000894 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000015c),
    .Q(sig00000194)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000895 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000179),
    .Q(sig0000015d),
    .Q15(NLW_blk00000895_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000896 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000015d),
    .Q(sig00000195)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000897 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000017a),
    .Q(sig0000015e),
    .Q15(NLW_blk00000897_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000898 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000015e),
    .Q(sig00000196)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000899 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000017b),
    .Q(sig0000015f),
    .Q15(NLW_blk00000899_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000089a (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000015f),
    .Q(sig00000197)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000089b (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000017e),
    .Q(sig00000162),
    .Q15(NLW_blk0000089b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000089c (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000162),
    .Q(sig0000019a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000089d (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000017c),
    .Q(sig00000160),
    .Q15(NLW_blk0000089d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000089e (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000160),
    .Q(sig00000198)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000089f (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000017d),
    .Q(sig00000161),
    .Q15(NLW_blk0000089f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008a0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000161),
    .Q(sig00000199)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008a1 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000180),
    .Q(sig00000164),
    .Q15(NLW_blk000008a1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008a2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000164),
    .Q(sig0000019c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008a3 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000181),
    .Q(sig00000165),
    .Q15(NLW_blk000008a3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008a4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000165),
    .Q(sig0000019d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008a5 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000182),
    .Q(sig00000166),
    .Q15(NLW_blk000008a5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008a6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000166),
    .Q(sig0000019e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008a7 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000183),
    .Q(sig00000167),
    .Q15(NLW_blk000008a7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008a8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000167),
    .Q(sig0000019f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008a9 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000184),
    .Q(sig00000168),
    .Q15(NLW_blk000008a9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008aa (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000168),
    .Q(sig000001a0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008ab (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000185),
    .Q(sig00000169),
    .Q15(NLW_blk000008ab_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008ac (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000169),
    .Q(sig000001a1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008ad (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001dd),
    .Q(sig000001ab),
    .Q15(NLW_blk000008ad_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008ae (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001ab),
    .Q(sig000001c4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008af (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000186),
    .Q(sig0000016a),
    .Q15(NLW_blk000008af_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008b0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000016a),
    .Q(sig000001a2)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008b1 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000187),
    .Q(sig0000016b),
    .Q15(NLW_blk000008b1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008b2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig0000016b),
    .Q(sig000001a3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008b3 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001de),
    .Q(sig000001ac),
    .Q15(NLW_blk000008b3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008b4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001ac),
    .Q(sig000001c5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008b5 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e9),
    .Q(sig000001b7),
    .Q15(NLW_blk000008b5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008b6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b7),
    .Q(sig000001d0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008b7 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001ef),
    .Q(sig000001bd),
    .Q15(NLW_blk000008b7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008b8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001bd),
    .Q(sig000001d6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008b9 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001f0),
    .Q(sig000001be),
    .Q15(NLW_blk000008b9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008ba (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001be),
    .Q(sig000001d7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008bb (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001f1),
    .Q(sig000001bf),
    .Q15(NLW_blk000008bb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008bc (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001bf),
    .Q(sig000001d8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008bd (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001f2),
    .Q(sig000001c0),
    .Q15(NLW_blk000008bd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008be (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001c0),
    .Q(sig000001d9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008bf (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001f5),
    .Q(sig000001c3),
    .Q15(NLW_blk000008bf_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008c0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001c3),
    .Q(sig000001dc)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008c1 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001f3),
    .Q(sig000001c1),
    .Q15(NLW_blk000008c1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008c2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001c1),
    .Q(sig000001da)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008c3 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001f4),
    .Q(sig000001c2),
    .Q15(NLW_blk000008c3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008c4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001c2),
    .Q(sig000001db)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008c5 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001df),
    .Q(sig000001ad),
    .Q15(NLW_blk000008c5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008c6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001ad),
    .Q(sig000001c6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008c7 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e0),
    .Q(sig000001ae),
    .Q15(NLW_blk000008c7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008c8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001ae),
    .Q(sig000001c7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008c9 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e3),
    .Q(sig000001b1),
    .Q15(NLW_blk000008c9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008ca (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b1),
    .Q(sig000001ca)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008cb (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e1),
    .Q(sig000001af),
    .Q15(NLW_blk000008cb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008cc (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001af),
    .Q(sig000001c8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008cd (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e2),
    .Q(sig000001b0),
    .Q15(NLW_blk000008cd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008ce (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b0),
    .Q(sig000001c9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008cf (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e4),
    .Q(sig000001b2),
    .Q15(NLW_blk000008cf_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008d0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b2),
    .Q(sig000001cb)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008d1 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e5),
    .Q(sig000001b3),
    .Q15(NLW_blk000008d1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008d2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b3),
    .Q(sig000001cc)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008d3 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e8),
    .Q(sig000001b6),
    .Q15(NLW_blk000008d3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008d4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b6),
    .Q(sig000001cf)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008d5 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e6),
    .Q(sig000001b4),
    .Q15(NLW_blk000008d5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008d6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b4),
    .Q(sig000001cd)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008d7 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001e7),
    .Q(sig000001b5),
    .Q15(NLW_blk000008d7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008d8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b5),
    .Q(sig000001ce)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008d9 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001ea),
    .Q(sig000001b8),
    .Q15(NLW_blk000008d9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008da (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b8),
    .Q(sig000001d1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008db (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001eb),
    .Q(sig000001b9),
    .Q15(NLW_blk000008db_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008dc (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001b9),
    .Q(sig000001d2)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008dd (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001ec),
    .Q(sig000001ba),
    .Q15(NLW_blk000008dd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008de (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001ba),
    .Q(sig000001d3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008df (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001ed),
    .Q(sig000001bb),
    .Q15(NLW_blk000008df_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008e0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001bb),
    .Q(sig000001d4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008e1 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000001ee),
    .Q(sig000001bc),
    .Q15(NLW_blk000008e1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008e2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000001bc),
    .Q(sig000001d5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008e3 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004ce),
    .Q(sig000004cd),
    .Q15(NLW_blk000008e3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008e4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004cd),
    .Q(sig000004cf)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008e5 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004df),
    .Q(sig000004db),
    .Q15(NLW_blk000008e5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008e6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004db),
    .Q(sig000004dd)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008e7 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000002b5),
    .Q(sig00000519),
    .Q15(NLW_blk000008e7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008e8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000519),
    .Q(sig0000051a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008e9 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004e0),
    .Q(sig000004dc),
    .Q15(NLW_blk000008e9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008ea (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004dc),
    .Q(sig000004de)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008eb (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004d9),
    .Q(sig000004d7),
    .Q15(NLW_blk000008eb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008ec (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004d7),
    .Q(sig000004d8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008ed (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004ad),
    .Q(sig000004b9),
    .Q15(NLW_blk000008ed_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008ee (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004b9),
    .Q(sig000004c4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008ef (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004b6),
    .Q(sig000004c1),
    .Q15(NLW_blk000008ef_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008f0 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004c1),
    .Q(sig000004cc)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008f1 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004b5),
    .Q(sig000004c0),
    .Q15(NLW_blk000008f1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008f2 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004c0),
    .Q(sig000004cb)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008f3 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004b4),
    .Q(sig000004bf),
    .Q15(NLW_blk000008f3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008f4 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004bf),
    .Q(sig000004ca)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008f5 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004b3),
    .Q(sig000004be),
    .Q15(NLW_blk000008f5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008f6 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004be),
    .Q(sig000004c9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008f7 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004b0),
    .Q(sig000004bb),
    .Q15(NLW_blk000008f7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008f8 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004bb),
    .Q(sig000004c6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008f9 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004b2),
    .Q(sig000004bd),
    .Q15(NLW_blk000008f9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008fa (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004bd),
    .Q(sig000004c8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008fb (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004b1),
    .Q(sig000004bc),
    .Q15(NLW_blk000008fb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008fc (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004bc),
    .Q(sig000004c7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008fd (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004af),
    .Q(sig000004ba),
    .Q15(NLW_blk000008fd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000008fe (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004ba),
    .Q(sig000004c5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000008ff (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004ac),
    .Q(sig000004b8),
    .Q15(NLW_blk000008ff_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000900 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004b8),
    .Q(sig000004c3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000901 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig000004ab),
    .Q(sig000004b7),
    .Q15(NLW_blk00000901_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000902 (
    .C(clk),
    .CE(sig00000002),
    .D(sig000004b7),
    .Q(sig000004c2)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000903 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000896),
    .Q(sig00000629),
    .Q15(NLW_blk00000903_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000904 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000629),
    .Q(sig0000062b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000905 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig00000897),
    .Q(sig00000628),
    .Q15(NLW_blk00000905_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000906 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000628),
    .Q(sig0000062a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000907 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(sig00000002),
    .CLK(clk),
    .D(sig0000035b),
    .Q(sig00000893),
    .Q15(NLW_blk00000907_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000908 (
    .C(clk),
    .CE(sig00000002),
    .D(sig00000893),
    .Q(sig00000894)
  );
// synthesis translate_on
endmodule