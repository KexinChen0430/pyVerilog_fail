module top ;
          wire  Net_432;
    electrical  Net_431;
          wire  Net_430;
          wire  Net_429;
          wire  Net_428;
    electrical  Net_427;
          wire  Net_345;
          wire  Net_344;
          wire  Net_343;
          wire  Net_342;
          wire  Net_341;
          wire  Net_340;
          wire  Net_338;
          wire  Net_337;
          wire  Net_336;
          wire  Net_335;
          wire  Net_333;
          wire  Net_339;
          wire  Net_334;
          wire  Net_291;
          wire  Net_290;
          wire  Net_289;
          wire  Net_288;
          wire  Net_433;
          wire  Net_293;
          wire  Net_212;
          wire  Net_211;
          wire  Net_210;
          wire  Net_208;
          wire  Net_207;
          wire  Net_206;
          wire  Net_204;
          wire  Net_203;
          wire  Net_202;
          wire  Net_201;
          wire  Net_200;
          wire  Net_199;
    electrical  Net_198;
    electrical  Net_197;
    electrical  Net_196;
    electrical  Net_195;
    electrical  Net_194;
    electrical  Net_193;
    electrical  Net_192;
    electrical  Net_191;
    electrical  Net_190;
    electrical  Net_189;
    electrical  Net_188;
    electrical  Net_187;
    electrical  Net_186;
    electrical  Net_185;
    electrical  Net_184;
    electrical  Net_183;
    electrical  Net_182;
    electrical  Net_181;
    electrical  Net_180;
    electrical  Net_179;
    electrical  Net_178;
    electrical  Net_177;
    electrical  Net_176;
    electrical  Net_175;
    electrical  Net_174;
    electrical  Net_173;
    electrical  Net_172;
    electrical  Net_171;
    electrical  Net_170;
    electrical  Net_169;
    electrical  Net_168;
    electrical  Net_167;
    electrical  Net_166;
    electrical  Net_165;
    electrical  Net_164;
    electrical  Net_163;
    electrical  Net_162;
    electrical  Net_161;
    electrical  Net_160;
    electrical  Net_159;
    electrical  Net_158;
    electrical  Net_157;
    electrical  Net_156;
    electrical  Net_155;
    electrical  Net_154;
    electrical  Net_153;
    electrical  Net_152;
    electrical  Net_151;
    electrical  Net_150;
    electrical  Net_149;
    electrical  Net_148;
    electrical  Net_147;
    electrical  Net_146;
    electrical  Net_145;
    electrical  Net_144;
    electrical  Net_143;
    electrical  Net_142;
    electrical  Net_141;
    electrical  Net_140;
    electrical  Net_139;
    electrical  Net_138;
    electrical  Net_137;
    electrical  Net_136;
    electrical  Net_135;
    electrical  Net_134;
    electrical  Net_133;
    electrical  Net_132;
    electrical  Net_131;
    electrical  Net_130;
    electrical  Net_129;
    electrical  Net_128;
    electrical  Net_127;
    electrical  Net_126;
    electrical  Net_125;
    electrical  Net_124;
    electrical  Net_123;
    electrical  Net_122;
    electrical  Net_121;
    electrical  Net_120;
    electrical  Net_119;
    electrical  Net_118;
    electrical  Net_117;
    electrical  Net_116;
    electrical  Net_115;
    electrical  Net_114;
    electrical  Net_113;
    electrical  Net_112;
    electrical  Net_111;
    electrical  Net_110;
    electrical  Net_109;
    electrical  Net_108;
    electrical  Net_107;
    electrical  Net_106;
    electrical  Net_105;
    electrical  Net_104;
    electrical  Net_103;
          wire  Net_102;
          wire  Net_101;
          wire  Net_100;
          wire  Net_99;
    electrical  Net_98;
    electrical  Net_97;
    electrical  Net_96;
    electrical  Net_95;
    electrical  Net_94;
    electrical  Net_93;
    electrical  Net_92;
    electrical  Net_91;
    electrical  Net_90;
    electrical  Net_89;
    electrical  Net_88;
    electrical  Net_87;
    electrical  Net_86;
    electrical  Net_85;
    electrical  Net_84;
    electrical  Net_83;
    electrical  Net_82;
    electrical  Net_81;
    electrical  Net_80;
    electrical  Net_79;
    electrical  Net_78;
    electrical  Net_77;
    electrical  Net_76;
    electrical  Net_75;
    electrical  Net_74;
    electrical  Net_73;
    electrical  Net_72;
    electrical  Net_71;
    electrical  Net_70;
    electrical  Net_69;
    electrical  Net_68;
    electrical  Net_67;
    electrical  Net_66;
    electrical  Net_65;
    electrical  Net_64;
    electrical  Net_63;
    electrical  Net_62;
    electrical  Net_61;
    electrical  Net_60;
    electrical  Net_59;
    electrical  Net_58;
    electrical  Net_57;
    electrical  Net_56;
    electrical  Net_55;
    electrical  Net_54;
    electrical  Net_53;
    electrical  Net_52;
    electrical  Net_51;
    electrical  Net_50;
    electrical  Net_49;
    electrical  Net_48;
    electrical  Net_47;
    electrical  Net_46;
    electrical  Net_45;
    electrical  Net_44;
    electrical  Net_43;
    electrical  Net_42;
    electrical  Net_41;
    electrical  Net_40;
    electrical  Net_39;
    electrical  Net_38;
    electrical  Net_37;
    electrical  Net_36;
    electrical  Net_35;
    electrical  Net_34;
    electrical  Net_33;
    electrical  Net_32;
    electrical  Net_31;
    electrical  Net_30;
    electrical  Net_29;
    electrical  Net_28;
    electrical  Net_27;
    electrical  Net_26;
    electrical  Net_25;
    electrical  Net_24;
    electrical  Net_23;
    electrical  Net_22;
    electrical  Net_21;
    electrical  Net_20;
    electrical  Net_19;
    electrical  Net_18;
    electrical  Net_17;
    electrical  Net_16;
    electrical  Net_15;
    electrical  Net_14;
    electrical  Net_13;
    electrical  Net_12;
    electrical  Net_11;
    electrical  Net_10;
    electrical  Net_9;
    electrical  Net_8;
    electrical  Net_7;
    electrical  Net_6;
    electrical  Net_5;
          wire  Net_4;
          wire  Net_3;
          wire  Net_2;
          wire  Net_1;
          wire  Net_205;
    electrical  Net_420;
          wire  Net_209;
          wire  Net_1822;
          wire  Net_286;
          wire  Net_284;
    electrical  Net_908;
    electrical  Net_907;
    ADC_SAR_SEQ_v2_0_1 TPS_ADC (
        .soc(1'b0),
        .aclk(1'b0),
        .sdone(Net_3),
        .eoc(Net_4),
        .AIN_10(Net_907),
        .AIN1(Net_908),
        .AIN_20(Net_5),
        .AIN_21(Net_6),
        .AIN_30(Net_7),
        .AIN_31(Net_8),
        .AIN3(Net_9),
        .AIN_40(Net_10),
        .AIN_41(Net_11),
        .AIN_50(Net_12),
        .AIN_51(Net_13),
        .AIN5(Net_14),
        .AIN_60(Net_15),
        .AIN_61(Net_16),
        .AIN_70(Net_17),
        .AIN_71(Net_18),
        .AIN7(Net_19),
        .AIN_80(Net_20),
        .AIN_81(Net_21),
        .AIN_90(Net_22),
        .AIN_91(Net_23),
        .AIN9(Net_24),
        .AIN_100(Net_25),
        .AIN_101(Net_26),
        .AIN_110(Net_27),
        .AIN_111(Net_28),
        .AIN11(Net_29),
        .AIN_120(Net_30),
        .AIN_121(Net_31),
        .AIN_130(Net_32),
        .AIN_131(Net_33),
        .AIN13(Net_34),
        .AIN_140(Net_35),
        .AIN_141(Net_36),
        .AIN_150(Net_37),
        .AIN_151(Net_38),
        .AIN15(Net_39),
        .AIN_160(Net_40),
        .AIN_161(Net_41),
        .AIN_170(Net_42),
        .AIN_171(Net_43),
        .AIN17(Net_44),
        .AIN_180(Net_45),
        .AIN_181(Net_46),
        .AIN_190(Net_47),
        .AIN_191(Net_48),
        .AIN19(Net_49),
        .AIN_200(Net_50),
        .AIN_201(Net_51),
        .AIN_210(Net_52),
        .AIN_211(Net_53),
        .AIN21(Net_54),
        .AIN_220(Net_55),
        .AIN_221(Net_56),
        .AIN_230(Net_57),
        .AIN_231(Net_58),
        .AIN23(Net_59),
        .AIN_240(Net_60),
        .AIN_241(Net_61),
        .AIN_250(Net_62),
        .AIN_251(Net_63),
        .AIN25(Net_64),
        .AIN_260(Net_65),
        .AIN_261(Net_66),
        .AIN_270(Net_67),
        .AIN_271(Net_68),
        .AIN27(Net_69),
        .AIN_280(Net_70),
        .AIN_281(Net_71),
        .AIN_290(Net_72),
        .AIN_291(Net_73),
        .AIN29(Net_74),
        .AIN_300(Net_75),
        .AIN_301(Net_76),
        .AIN_310(Net_77),
        .AIN_311(Net_78),
        .AIN31(Net_79),
        .AIN_320(Net_80),
        .AIN_321(Net_81),
        .AIN49(Net_82),
        .AIN50(Net_83),
        .AIN51(Net_84),
        .AIN52(Net_85),
        .AIN53(Net_86),
        .AIN54(Net_87),
        .AIN55(Net_88),
        .AIN56(Net_89),
        .AIN57(Net_90),
        .AIN58(Net_91),
        .AIN59(Net_92),
        .AIN60(Net_93),
        .AIN61(Net_94),
        .AIN62(Net_95),
        .AIN63(Net_96),
        .AIN64(Net_97),
        .vdac_ref(Net_98));
	wire [0:0] tmpOE__TPS_0_net;
	wire [0:0] tmpFB_0__TPS_0_net;
	wire [0:0] tmpIO_0__TPS_0_net;
	wire [0:0] tmpINTERRUPT_0__TPS_0_net;
	electrical [0:0] tmpSIOVREF__TPS_0_net;
	cy_psoc3_pins_v1_10
		#(.id("77715107-f8d5-47e5-a629-0fb83101ac6b"),
		  .drive_mode(3'b011),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("A"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		TPS_0
		 (.oe(tmpOE__TPS_0_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__TPS_0_net[0:0]}),
		  .analog({Net_907}),
		  .io({tmpIO_0__TPS_0_net[0:0]}),
		  .siovref(tmpSIOVREF__TPS_0_net),
		  .interrupt({tmpINTERRUPT_0__TPS_0_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__TPS_0_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__TPS_1_net;
	wire [0:0] tmpFB_0__TPS_1_net;
	wire [0:0] tmpIO_0__TPS_1_net;
	wire [0:0] tmpINTERRUPT_0__TPS_1_net;
	electrical [0:0] tmpSIOVREF__TPS_1_net;
	cy_psoc3_pins_v1_10
		#(.id("14425a1b-440b-4507-9dac-74192c9da648"),
		  .drive_mode(3'b011),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("A"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		TPS_1
		 (.oe(tmpOE__TPS_1_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__TPS_1_net[0:0]}),
		  .analog({Net_908}),
		  .io({tmpIO_0__TPS_1_net[0:0]}),
		  .siovref(tmpSIOVREF__TPS_1_net),
		  .interrupt({tmpINTERRUPT_0__TPS_1_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__TPS_1_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    ADC_SAR_SEQ_v2_0_3 APPS_ADC (
        .soc(1'b0),
        .aclk(1'b0),
        .sdone(Net_101),
        .eoc(Net_102),
        .AIN_10(Net_103),
        .AIN1(Net_104),
        .AIN_20(Net_105),
        .AIN_21(Net_106),
        .AIN_30(Net_107),
        .AIN_31(Net_108),
        .AIN3(Net_109),
        .AIN_40(Net_110),
        .AIN_41(Net_111),
        .AIN_50(Net_112),
        .AIN_51(Net_113),
        .AIN5(Net_114),
        .AIN_60(Net_115),
        .AIN_61(Net_116),
        .AIN_70(Net_117),
        .AIN_71(Net_118),
        .AIN7(Net_119),
        .AIN_80(Net_120),
        .AIN_81(Net_121),
        .AIN_90(Net_122),
        .AIN_91(Net_123),
        .AIN9(Net_124),
        .AIN_100(Net_125),
        .AIN_101(Net_126),
        .AIN_110(Net_127),
        .AIN_111(Net_128),
        .AIN11(Net_129),
        .AIN_120(Net_130),
        .AIN_121(Net_131),
        .AIN_130(Net_132),
        .AIN_131(Net_133),
        .AIN13(Net_134),
        .AIN_140(Net_135),
        .AIN_141(Net_136),
        .AIN_150(Net_137),
        .AIN_151(Net_138),
        .AIN15(Net_139),
        .AIN_160(Net_140),
        .AIN_161(Net_141),
        .AIN_170(Net_142),
        .AIN_171(Net_143),
        .AIN17(Net_144),
        .AIN_180(Net_145),
        .AIN_181(Net_146),
        .AIN_190(Net_147),
        .AIN_191(Net_148),
        .AIN19(Net_149),
        .AIN_200(Net_150),
        .AIN_201(Net_151),
        .AIN_210(Net_152),
        .AIN_211(Net_153),
        .AIN21(Net_154),
        .AIN_220(Net_155),
        .AIN_221(Net_156),
        .AIN_230(Net_157),
        .AIN_231(Net_158),
        .AIN23(Net_159),
        .AIN_240(Net_160),
        .AIN_241(Net_161),
        .AIN_250(Net_162),
        .AIN_251(Net_163),
        .AIN25(Net_164),
        .AIN_260(Net_165),
        .AIN_261(Net_166),
        .AIN_270(Net_167),
        .AIN_271(Net_168),
        .AIN27(Net_169),
        .AIN_280(Net_170),
        .AIN_281(Net_171),
        .AIN_290(Net_172),
        .AIN_291(Net_173),
        .AIN29(Net_174),
        .AIN_300(Net_175),
        .AIN_301(Net_176),
        .AIN_310(Net_177),
        .AIN_311(Net_178),
        .AIN31(Net_179),
        .AIN_320(Net_180),
        .AIN_321(Net_181),
        .AIN49(Net_182),
        .AIN50(Net_183),
        .AIN51(Net_184),
        .AIN52(Net_185),
        .AIN53(Net_186),
        .AIN54(Net_187),
        .AIN55(Net_188),
        .AIN56(Net_189),
        .AIN57(Net_190),
        .AIN58(Net_191),
        .AIN59(Net_192),
        .AIN60(Net_193),
        .AIN61(Net_194),
        .AIN62(Net_195),
        .AIN63(Net_196),
        .AIN64(Net_197),
        .vdac_ref(Net_198));
	wire [0:0] tmpOE__APPS_0_net;
	wire [0:0] tmpFB_0__APPS_0_net;
	wire [0:0] tmpIO_0__APPS_0_net;
	wire [0:0] tmpINTERRUPT_0__APPS_0_net;
	electrical [0:0] tmpSIOVREF__APPS_0_net;
	cy_psoc3_pins_v1_10
		#(.id("6508d192-65fb-4cff-b19b-01459585c961"),
		  .drive_mode(3'b011),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("A"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		APPS_0
		 (.oe(tmpOE__APPS_0_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__APPS_0_net[0:0]}),
		  .analog({Net_103}),
		  .io({tmpIO_0__APPS_0_net[0:0]}),
		  .siovref(tmpSIOVREF__APPS_0_net),
		  .interrupt({tmpINTERRUPT_0__APPS_0_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__APPS_0_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__APPS_1_net;
	wire [0:0] tmpFB_0__APPS_1_net;
	wire [0:0] tmpIO_0__APPS_1_net;
	wire [0:0] tmpINTERRUPT_0__APPS_1_net;
	electrical [0:0] tmpSIOVREF__APPS_1_net;
	cy_psoc3_pins_v1_10
		#(.id("5e195aa5-59f6-4b8b-b29d-3cc2166d48ca"),
		  .drive_mode(3'b011),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("A"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		APPS_1
		 (.oe(tmpOE__APPS_1_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__APPS_1_net[0:0]}),
		  .analog({Net_104}),
		  .io({tmpIO_0__APPS_1_net[0:0]}),
		  .siovref(tmpSIOVREF__APPS_1_net),
		  .interrupt({tmpINTERRUPT_0__APPS_1_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__APPS_1_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    PWM_v3_30_4 SERVO_PWM (
        .reset(1'b0),
        .clock(Net_1822),
        .tc(Net_200),
        .pwm1(Net_201),
        .pwm2(Net_202),
        .interrupt(Net_203),
        .capture(1'b0),
        .kill(Net_205),
        .enable(1'b1),
        .trigger(1'b0),
        .cmp_sel(1'b0),
        .pwm(Net_209),
        .ph1(Net_210),
        .ph2(Net_211));
    defparam SERVO_PWM.Resolution = 16;
	wire [0:0] tmpOE__SERVO_OUT_net;
	wire [0:0] tmpFB_0__SERVO_OUT_net;
	wire [0:0] tmpIO_0__SERVO_OUT_net;
	wire [0:0] tmpINTERRUPT_0__SERVO_OUT_net;
	electrical [0:0] tmpSIOVREF__SERVO_OUT_net;
	cy_psoc3_pins_v1_10
		#(.id("e851a3b9-efb8-48be-bbb8-b303b216c393"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		SERVO_OUT
		 (.oe(tmpOE__SERVO_OUT_net),
		  .y({Net_209}),
		  .fb({tmpFB_0__SERVO_OUT_net[0:0]}),
		  .io({tmpIO_0__SERVO_OUT_net[0:0]}),
		  .siovref(tmpSIOVREF__SERVO_OUT_net),
		  .interrupt({tmpINTERRUPT_0__SERVO_OUT_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__SERVO_OUT_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	cy_clock_v1_0
		#(.id("8d232960-f3fa-479f-8ed8-8a4839b5bc1f"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("1000000000"),
		  .is_direct(0),
		  .is_digital(1))
		pwm_clock
		 (.clock_out(Net_1822));
	cy_clock_v1_0
		#(.id("c0fb34bd-1044-4931-9788-16b01ce89812"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("31250000000"),
		  .is_direct(0),
		  .is_digital(1))
		timer_clock
		 (.clock_out(Net_284));
    ZeroTerminal ZeroTerminal_1 (
        .z(Net_286));
    Timer_v2_70_5 Timer (
        .reset(Net_286),
        .interrupt(Net_433),
        .enable(1'b1),
        .trigger(1'b1),
        .capture(1'b0),
        .capture_out(Net_291),
        .tc(Net_205),
        .clock(Net_284));
    defparam Timer.CaptureCount = 2;
    defparam Timer.CaptureCounterEnabled = 0;
    defparam Timer.DeviceFamily = "PSoC5";
    defparam Timer.InterruptOnCapture = 0;
    defparam Timer.InterruptOnTC = 1;
    defparam Timer.Resolution = 16;
    defparam Timer.SiliconRevision = "0";
	wire [0:0] tmpOE__Tx_1_net;
	wire [0:0] tmpFB_0__Tx_1_net;
	wire [0:0] tmpIO_0__Tx_1_net;
	wire [0:0] tmpINTERRUPT_0__Tx_1_net;
	electrical [0:0] tmpSIOVREF__Tx_1_net;
	cy_psoc3_pins_v1_10
		#(.id("ed092b9b-d398-4703-be89-cebf998501f6"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		Tx_1
		 (.oe(tmpOE__Tx_1_net),
		  .y({Net_334}),
		  .fb({tmpFB_0__Tx_1_net[0:0]}),
		  .io({tmpIO_0__Tx_1_net[0:0]}),
		  .siovref(tmpSIOVREF__Tx_1_net),
		  .interrupt({tmpINTERRUPT_0__Tx_1_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__Tx_1_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__Rx_1_net;
	wire [0:0] tmpIO_0__Rx_1_net;
	wire [0:0] tmpINTERRUPT_0__Rx_1_net;
	electrical [0:0] tmpSIOVREF__Rx_1_net;
	cy_psoc3_pins_v1_10
		#(.id("1425177d-0d0e-4468-8bcc-e638e5509a9b"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		Rx_1
		 (.oe(tmpOE__Rx_1_net),
		  .y({1'b0}),
		  .fb({Net_339}),
		  .io({tmpIO_0__Rx_1_net[0:0]}),
		  .siovref(tmpSIOVREF__Rx_1_net),
		  .interrupt({tmpINTERRUPT_0__Rx_1_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__Rx_1_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    UART_v2_50_6 UART (
        .cts_n(1'b0),
        .tx(Net_334),
        .rts_n(Net_335),
        .tx_en(Net_336),
        .clock(1'b0),
        .reset(1'b0),
        .rx(Net_339),
        .tx_interrupt(Net_340),
        .rx_interrupt(Net_341),
        .tx_data(Net_342),
        .tx_clk(Net_343),
        .rx_data(Net_344),
        .rx_clk(Net_345));
    defparam UART.Address1 = 0;
    defparam UART.Address2 = 0;
    defparam UART.EnIntRXInterrupt = 0;
    defparam UART.EnIntTXInterrupt = 0;
    defparam UART.FlowControl = 0;
    defparam UART.HalfDuplexEn = 0;
    defparam UART.HwTXEnSignal = 1;
    defparam UART.NumDataBits = 8;
    defparam UART.NumStopBits = 1;
    defparam UART.ParityType = 0;
    defparam UART.RXEnable = 1;
    defparam UART.TXEnable = 1;
    ADC_DelSig_v3_20_7 BRAKE_ADC (
        .vplus(Net_420),
        .vminus(Net_427),
        .soc(1'b1),
        .eoc(Net_429),
        .aclk(1'b0),
        .nVref(Net_431),
        .mi(1'b0));
	wire [0:0] tmpOE__BRAKE_net;
	wire [0:0] tmpFB_0__BRAKE_net;
	wire [0:0] tmpIO_0__BRAKE_net;
	wire [0:0] tmpINTERRUPT_0__BRAKE_net;
	electrical [0:0] tmpSIOVREF__BRAKE_net;
	cy_psoc3_pins_v1_10
		#(.id("029dc6f8-8ce0-418b-bd71-68702303c56b"),
		  .drive_mode(3'b000),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("A"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		BRAKE
		 (.oe(tmpOE__BRAKE_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__BRAKE_net[0:0]}),
		  .analog({Net_420}),
		  .io({tmpIO_0__BRAKE_net[0:0]}),
		  .siovref(tmpSIOVREF__BRAKE_net),
		  .interrupt({tmpINTERRUPT_0__BRAKE_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__BRAKE_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
endmodule