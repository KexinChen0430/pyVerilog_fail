module bug778 ();
   virtual if_bug777.master bar;
endmodule