module  xye129(
   sys_clk,
   rst_n,
   dmfe774,
   hb7e87f,
   al4bbdd,
   qgcbe8c,
   fn5f460,
   ayfa306,
   sj397d1,
   thec436,
   ui621b7,
   uk10db8,
   ng86dc0,
   cb36e02,
   pub7014,
   twb80a3,
   zkc051a,
   ux28d2,
   fc14694,
   aaa34a3,
   qi1a518,
   nrd28c0,
   ph94607,
   coa303f,
   ir181f8,
   dmc0fc5
   );
parameter ep7e2b    = 3'b000;
parameter hq3f15c   = 3'b001;
parameter mrf8ae3  = 3'b010;
parameter zkc571d    = 3'b011;
parameter sw2b8ea   = 3'b100;
parameter me5c751  = 3'b101;
parameter uvc3724   = 2'b00;
parameter je1b925  = 2'b01;
parameter mrdc92b = 2'b10;
input                     sys_clk;
input                     rst_n;
input                     dmfe774;
input                     hb7e87f;
input  [2:0]              al4bbdd;
input                     qgcbe8c;
input                     fn5f460;
input                     ayfa306;
input  [1:0]              sj397d1;
input  [2:0]              thec436;
input  [19:0]             ui621b7;
input                     uk10db8;
input                     ng86dc0;
input                     cb36e02;
input  [15:0]             pub7014;
input                     twb80a3;
input                     zkc051a;
input                     ux28d2;
input                     fc14694;
output                    aaa34a3;
output  [8:0]             qi1a518;
output  [12:0]            nrd28c0;
output  [8:0]             ph94607;
output  [12:0]            coa303f;
output  [8:0]             ir181f8;
output  [12:0]            dmc0fc5;
reg     [8:0]             qi1a518;
reg     [12:0]            nrd28c0;
reg     [8:0]             ph94607;
reg     [12:0]            coa303f;
reg     [8:0]             ir181f8;
reg     [12:0]            dmc0fc5;
reg  [11:0]               hb7edba;
reg  [7:0]                jpf6dd6;
reg                       ri11ac4;
reg                       ale2358;
reg  [11:0]               fpbad83;
reg  [7:0]                shd6c1e;
reg                       pf6b110;
reg                       ou8d622;
reg  [11:0]               ng83d4e;
reg  [7:0]                ba1ea72;
reg                       wwc4432;
reg                       lq58886;
reg                       ip4e4c0;
reg                       ui72605;
reg                       hq93029;
reg  [11:0]               mg9814a;
reg  [7:0]                jcc0a51;
reg  [11:0]               ym528b;
reg  [7:0]                mt29458;
reg  [11:0]               th4a2c5;
reg  [7:0]                gb5162f;
reg                       lf8b17d;
reg                       tu58bef;
reg                       jcc5f7a;
reg                       zm2fbd3;
reg  [8:0]                qg7de9b;
reg                       eaef4d9;
reg                       cz7a6c8;
reg                       yxd3645;
reg                       vx9b22c;
reg                       ald9166;
reg                       thc8b35;
reg                       hb459af;
reg                       kf2cd7f;
reg                       xw66bfc;
reg                       xy35fe3;
reg                       hdaff1b;
reg                       en7f8df;
reg                       ldfc6fc;
reg                       pfe37e6;
reg  [11:0]               hq1bf36;
reg  [7:0]                vidf9b3;
reg  [11:0]               fnfcd9b;
reg  [7:0]                xje6cdf;
reg                       yz366ff;
reg                       mgb37fd;
reg                       xl9bfe9;
reg                       tudff4f;
reg                       meffa7b;
reg                       wjfd3d8;
reg [1:0]                 zxe9ec4;
reg [4:0]                 pf4f626;
wire                      bl7b137;
wire                      rtd89bf;
wire [11:0]               suc4dfe;
wire [7:0]                ux26ff1;
wire                      bn37f8d;
wire                      jrbfc6e;
wire                      xwfe376;
wire                      jcf1bb3;
reg wy8dd9b;
reg alc3f66;
reg [2 : 0] ne766cf;
reg kf2c072;
reg cz60395;
reg ls1cad;
reg [1 : 0] pue56b;
reg [2 : 0] ld7b3a3;
reg [19 : 0] shd9d1f;
reg ayce8fc;
reg hb747e0;
reg coa3f06;
reg [15 : 0] ks1f831;
reg vvfc189;
reg ose0c4e;
reg bn6270;
reg mg31387;
reg [11 : 0] ri89c38;
reg [7 : 0] qt4e1c3;
reg ou8887d;
reg kd5110f;
reg [11 : 0] ph38769;
reg [7 : 0] uvc3b4e;
reg ou21f4c;
reg sh443e9;
reg [11 : 0] by69d25;
reg [7 : 0] en4e92a;
reg os7d300;
reg ymfa60;
reg xy2553c;
reg xy2a9e3;
reg cz54f1b;
reg [11 : 0] zma78dc;
reg [7 : 0] oh3c6e3;
reg [11 : 0] nre371c;
reg [7 : 0] ri1b8e6;
reg [11 : 0] yxdc733;
reg [7 : 0] dze399d;
reg vx1ccef;
reg ble677e;
reg an33bf6;
reg ym9dfb4;
reg [8 : 0] wwefda0;
reg vv7ed01;
reg rtf680e;
reg gdb4076;
reg xla03b4;
reg xy1da7;
reg hqed3b;
reg jc769da;
reg uxb4ed2;
reg hqa7695;
reg uk3b4aa;
reg lqda551;
reg zxd2a8a;
reg gd95457;
reg lfaa2bd;
reg [11 : 0] gb515ee;
reg [7 : 0] kf8af75;
reg [11 : 0] ho57bac;
reg [7 : 0] ribdd63;
reg neeeb1b;
reg al758db;
reg coac6dd;
reg ps636e9;
reg hq1b74a;
reg qgdba52;
reg [1 : 0] rtdd291;
reg [4 : 0] zxe948f;
reg th4a47f;
reg fa523ff;
reg [11 : 0] zz91ffa;
reg [7 : 0] cb8ffd6;
reg wj7feb4;
reg wwff5a4;
reg ayfad21;
reg end6908;
reg [2047:0] necf6c2;
wire [76:0] ld7b613;
localparam qgdb09f = 77,nrd84f8 = 32'hfdfff10b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
assign aaa34a3 = gd95457 | lfaa2bd;
assign suc4dfe = shd9d1f[11:0];
assign ux26ff1  = shd9d1f[19:12];
always @ (*) begin   hq1bf36 = 0;   vidf9b3  = 0;   case(pue56b)      uvc3724   : begin         hq1bf36 = ri89c38;         vidf9b3  = qt4e1c3;      end      je1b925  :  begin         hq1bf36 = ph38769;         vidf9b3  = uvc3b4e;      end      mrdc92b :  begin         hq1bf36 = by69d25;         vidf9b3  = en4e92a;      end   endcase
end
assign bn37f8d  = (cb8ffd6 != 0) ? 1'b1 : 1'b0;
assign jrbfc6e = (zz91ffa != 0) ? 1'b1 : 1'b0;
assign jcf1bb3 = neeeb1b | coac6dd | hq1b74a;
assign xwfe376  = al758db | ps636e9 | qgdba52;
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      ldfc6fc  <= 1'b0;      pfe37e6  <= 1'b0;      fnfcd9b         <= 0;      xje6cdf          <= 0;      yz366ff            <= 1'b0;      mgb37fd            <= 1'b0;      xl9bfe9           <= 1'b0;      tudff4f           <= 1'b0;      meffa7b          <= 1'b0;      wjfd3d8          <= 1'b0;   end   else begin      ldfc6fc  <= 1'b0;      pfe37e6  <= 1'b0;      yz366ff            <= 1'b0;      mgb37fd            <= 1'b0;      xl9bfe9           <= 1'b0;      tudff4f           <= 1'b0;      meffa7b          <= 1'b0;      wjfd3d8          <= 1'b0;            if(ld7b3a3 == ne766cf) begin         case(pue56b)            uvc3724 : begin               if(ls1cad && xy2553c) begin                  yz366ff <= !ou8887d;                  mgb37fd <= !kd5110f;                  if((ou8887d && wwff5a4) || (kd5110f && wj7feb4))                     ldfc6fc  <= 1'b1;               end            end            je1b925 : begin               if(ls1cad && xy2a9e3) begin                  xl9bfe9 <= !ou21f4c;                  tudff4f <= !sh443e9;                  if((ou21f4c && wwff5a4) || (sh443e9 && wj7feb4))                     ldfc6fc  <= 1'b1;               end            end            mrdc92b : begin               if(ls1cad && cz54f1b) begin                  meffa7b <= !os7d300;                  wjfd3d8 <= !ymfa60;                  if((os7d300 && wwff5a4) || (ymfa60 && wj7feb4))                     ldfc6fc  <= 1'b1;               end            end         endcase      end            fnfcd9b <= zz91ffa - gb515ee;      xje6cdf  <= cb8ffd6  - kf8af75;      if(((ho57bac > 2047) && end6908) || ((ribdd63 > 127) && ayfad21))         pfe37e6  <= 1'b1;      else         pfe37e6  <= 1'b0;   end
end
assign bl7b137  = kf2c072 | cz60395 | ls1cad;
assign rtd89bf     = kf2c072 | cz60395;
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      hb7edba      <= 12'h000;      jpf6dd6       <= 8'h00;      fpbad83     <= 12'h000;      shd6c1e      <= 8'h00;      ng83d4e    <= 12'h000;      ba1ea72     <= 8'h00;      ri11ac4        <= 1'b0;      ale2358        <= 1'b0;      pf6b110       <= 1'b0;      ou8d622       <= 1'b0;      wwc4432      <= 1'b0;      lq58886      <= 1'b0;      ip4e4c0          <= 1'b0;      ui72605         <= 1'b0;      hq93029        <= 1'b0;   end   else begin                                    if(ld7b3a3 == ne766cf) begin         case(pue56b)            uvc3724 : begin               if(th4a47f) begin                  hb7edba    <= zz91ffa;                  jpf6dd6     <= cb8ffd6;               end               if(fa523ff) begin                  if(xy2553c == 1'b0) begin                     ri11ac4      <= (wwff5a4) ? 1'b0 : 1'b1;                     ale2358      <= (wj7feb4) ? 1'b0 : 1'b1;                  end               end            end            je1b925 : begin               if(th4a47f) begin                  fpbad83   <= zz91ffa;                  shd6c1e    <= cb8ffd6;               end               if(fa523ff) begin                  if(xy2a9e3 == 1'b0) begin                     pf6b110     <= (wwff5a4) ? 1'b0 : 1'b1;                     ou8d622     <= (wj7feb4) ? 1'b0 : 1'b1;                  end               end            end            mrdc92b : begin               if(th4a47f) begin                  ng83d4e  <= zz91ffa;                  ba1ea72   <= cb8ffd6;               end               if(fa523ff) begin                  if(cz54f1b == 1'b0) begin                     wwc4432    <= (wwff5a4) ? 1'b0 : 1'b1;                     lq58886    <= (wj7feb4) ? 1'b0 : 1'b1;                  end               end            end         endcase      end                        if(wy8dd9b || !alc3f66) begin         ip4e4c0   <= 1'b0;         ui72605  <= 1'b0;         hq93029 <= 1'b0;      end      else if((ld7b3a3 == ne766cf) && fa523ff) begin         case(pue56b)            uvc3724   : ip4e4c0   <= 1'b1;            je1b925  : ui72605  <= 1'b1;            mrdc92b : hq93029 <= 1'b1;         endcase      end   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      lf8b17d     <= 1'b0;      zm2fbd3      <= 1'b0;      tu58bef  <= 1'b0;      jcc5f7a  <= 1'b0;   end   else begin      lf8b17d     <= ayce8fc;      zm2fbd3      <= coa3f06;      tu58bef  <= vx1ccef | bn6270 | vvfc189;      jcc5f7a  <= bn6270 | vvfc189;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      zxe9ec4   <= 2'b00;      pf4f626  <= 5'b00000;   end   else if (ayce8fc) begin      zxe9ec4   <= ks1f831[14:13];      pf4f626  <= ks1f831[12:8];   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      eaef4d9     <= 1'b0 ;      cz7a6c8     <= 1'b0 ;      yxd3645    <= 1'b0 ;      vx9b22c    <= 1'b0 ;      ald9166   <= 1'b0;      thc8b35   <= 1'b0;      qg7de9b <= 9'h000;      hb459af   <= 1'b0 ;      kf2cd7f   <= 1'b0 ;      xw66bfc  <= 1'b0 ;      xy35fe3  <= 1'b0 ;      hdaff1b <= 1'b0;      en7f8df <= 1'b0;   end   else begin                  if(mg31387 || ose0c4e)         qg7de9b <= 9'h001;      else if(vx1ccef) begin         if(ks1f831[1:0] == 2'b00)               qg7de9b <= {(~(|ks1f831[9:2])), ks1f831[9:2]};         else              qg7de9b <= ks1f831[9:2] + 1;      end      if(bn6270 || vvfc189) begin         if(bn6270) begin              if(!ymfa60)               ald9166 <= 1'b1;            if(!os7d300)               thc8b35 <= mg31387;         end         else begin              if(!kd5110f)               eaef4d9 <= 1'b1;            if(!ou8887d)               cz7a6c8 <= ose0c4e;         end      end      else if(vx1ccef) begin         if(!ou8887d)            cz7a6c8   <= (((zxe948f[4:3] == 2'b10) || (zxe948f[2:0] == 3'b000)) && rtdd291[1]) ? 1'b1 : 1'b0;         if(!kd5110f)            eaef4d9   <= ((zxe948f[4:3] == 2'b10) || ((zxe948f[2:0] == 3'b000) && rtdd291[1])) ? 1'b1 : 1'b0;         if(!ou21f4c)            vx9b22c  <= ((zxe948f[4:3] == 2'b00) && rtdd291[1] && (zxe948f[2:0] != 3'b000)) ? 1'b1 : 1'b0;         if(!sh443e9)            yxd3645  <= ((zxe948f[4:3] == 2'b00) && !((zxe948f[2:0] == 3'b000) && rtdd291[1])) ? 1'b1 : 1'b0;         if(!ymfa60)            ald9166 <= (zxe948f == 5'b0_1010) ? 1'b1 : 1'b0;         if(!os7d300)            thc8b35 <= ((zxe948f == 5'b0_1010) && rtdd291[1]) ? 1'b1 : 1'b0;      end      else if (hb747e0 || coa3f06 || an33bf6) begin         eaef4d9   <= 1'b0;         cz7a6c8   <= 1'b0;         yxd3645  <= 1'b0;         vx9b22c  <= 1'b0;         ald9166 <= 1'b0;         thc8b35 <= 1'b0;      end      hb459af   <= vv7ed01;      kf2cd7f   <= rtf680e;      xw66bfc  <= gdb4076;      xy35fe3  <= xla03b4;      hdaff1b <= xy1da7;      en7f8df <= hqed3b;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      jcc0a51    <= 8'h00;      mt29458   <= 8'h00;      gb5162f  <= 8'h00;      mg9814a   <= 12'h000;      th4a2c5 <= 12'h000;      ym528b  <= 12'h000;   end   else begin      if(wy8dd9b || !alc3f66) begin         jcc0a51    <= 8'h00;         mt29458   <= 8'h00;         gb5162f  <= 8'h00;         mg9814a   <= 12'h000;         th4a2c5 <= 12'h000;         ym528b  <= 12'h000;      end      else if(ble677e) begin         jcc0a51   <= (vv7ed01) ? (oh3c6e3 + 1'b1) : oh3c6e3;         mt29458  <= (gdb4076) ? (ri1b8e6 + 1'b1) : ri1b8e6;         gb5162f <= (xy1da7) ? (dze399d + 1'b1) : dze399d;         mg9814a   <= (rtf680e) ? (zma78dc + wwefda0) : zma78dc;         ym528b  <= (xla03b4) ? (nre371c + 1'b1) : nre371c;         th4a2c5 <= (hqed3b) ? (yxdc733 + wwefda0) : yxdc733;      end      else if(ym9dfb4) begin         jcc0a51   <= (jc769da) ? (oh3c6e3 - 1'b1) : oh3c6e3;         mt29458  <= (hqa7695) ? (ri1b8e6 - 1'b1) : ri1b8e6;         gb5162f <= (lqda551) ? (dze399d - 1'b1) : dze399d;         mg9814a   <= (uxb4ed2) ? (zma78dc - wwefda0) : zma78dc;         ym528b  <= (uk3b4aa) ? (nre371c - 1'b1) : nre371c;         th4a2c5 <= (zxd2a8a) ? (yxdc733 - wwefda0) : yxdc733;      end   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      qi1a518    <= 9'h00;      ph94607   <= 9'h00;      ir181f8  <= 9'h00;      nrd28c0    <= 13'h000;      coa303f   <= 13'h000;      dmc0fc5  <= 13'h000;   end   else begin      qi1a518[7:0]    <= qt4e1c3 - oh3c6e3;      ph94607[7:0]   <= uvc3b4e - ri1b8e6;      ir181f8[7:0]  <= en4e92a - dze399d;
      nrd28c0[11:0]   <= ri89c38 - zma78dc;      coa303f[11:0]  <= ph38769 - nre371c;      dmc0fc5[11:0] <= by69d25 - yxdc733;            qi1a518[8]      <= kd5110f;      ph94607[8]     <= sh443e9;      ir181f8[8]    <= ymfa60;      nrd28c0[12]     <= ou8887d;      coa303f[12]    <= ou21f4c;      dmc0fc5[12]   <= os7d300;   end
end
always@* begin wy8dd9b<=ld7b613[0];alc3f66<=ld7b613[1];ne766cf<={al4bbdd>>1,ld7b613[2]};kf2c072<=ld7b613[3];cz60395<=ld7b613[4];ls1cad<=ld7b613[5];pue56b<={sj397d1>>1,ld7b613[6]};ld7b3a3<={thec436>>1,ld7b613[7]};shd9d1f<={ui621b7>>1,ld7b613[8]};ayce8fc<=ld7b613[9];hb747e0<=ld7b613[10];coa3f06<=ld7b613[11];ks1f831<={pub7014>>1,ld7b613[12]};vvfc189<=ld7b613[13];ose0c4e<=ld7b613[14];bn6270<=ld7b613[15];mg31387<=ld7b613[16];ri89c38<={hb7edba>>1,ld7b613[17]};qt4e1c3<={jpf6dd6>>1,ld7b613[18]};ou8887d<=ld7b613[19];kd5110f<=ld7b613[20];ph38769<={fpbad83>>1,ld7b613[21]};uvc3b4e<={shd6c1e>>1,ld7b613[22]};ou21f4c<=ld7b613[23];sh443e9<=ld7b613[24];by69d25<={ng83d4e>>1,ld7b613[25]};en4e92a<={ba1ea72>>1,ld7b613[26]};os7d300<=ld7b613[27];ymfa60<=ld7b613[28];xy2553c<=ld7b613[29];xy2a9e3<=ld7b613[30];cz54f1b<=ld7b613[31];zma78dc<={mg9814a>>1,ld7b613[32]};oh3c6e3<={jcc0a51>>1,ld7b613[33]};nre371c<={ym528b>>1,ld7b613[34]};ri1b8e6<={mt29458>>1,ld7b613[35]};yxdc733<={th4a2c5>>1,ld7b613[36]};dze399d<={gb5162f>>1,ld7b613[37]};vx1ccef<=ld7b613[38];ble677e<=ld7b613[39];an33bf6<=ld7b613[40];ym9dfb4<=ld7b613[41];wwefda0<={qg7de9b>>1,ld7b613[42]};vv7ed01<=ld7b613[43];rtf680e<=ld7b613[44];gdb4076<=ld7b613[45];xla03b4<=ld7b613[46];xy1da7<=ld7b613[47];hqed3b<=ld7b613[48];jc769da<=ld7b613[49];uxb4ed2<=ld7b613[50];hqa7695<=ld7b613[51];uk3b4aa<=ld7b613[52];lqda551<=ld7b613[53];zxd2a8a<=ld7b613[54];gd95457<=ld7b613[55];lfaa2bd<=ld7b613[56];gb515ee<={hq1bf36>>1,ld7b613[57]};kf8af75<={vidf9b3>>1,ld7b613[58]};ho57bac<={fnfcd9b>>1,ld7b613[59]};ribdd63<={xje6cdf>>1,ld7b613[60]};neeeb1b<=ld7b613[61];al758db<=ld7b613[62];coac6dd<=ld7b613[63];ps636e9<=ld7b613[64];hq1b74a<=ld7b613[65];qgdba52<=ld7b613[66];rtdd291<={zxe9ec4>>1,ld7b613[67]};zxe948f<={pf4f626>>1,ld7b613[68]};th4a47f<=ld7b613[69];fa523ff<=ld7b613[70];zz91ffa<={suc4dfe>>1,ld7b613[71]};cb8ffd6<={ux26ff1>>1,ld7b613[72]};wj7feb4<=ld7b613[73];wwff5a4<=ld7b613[74];ayfad21<=ld7b613[75];end6908<=ld7b613[76];end
always@* begin necf6c2[2047]<=hb7e87f;necf6c2[2046]<=al4bbdd[0];necf6c2[2044]<=qgcbe8c;necf6c2[2040]<=fn5f460;necf6c2[2032]<=ayfa306;necf6c2[2016]<=sj397d1[0];necf6c2[1985]<=thec436[0];necf6c2[1950]<=hb7edba[0];necf6c2[1930]<=pf6b110;necf6c2[1923]<=ui621b7[0];necf6c2[1878]<=pfe37e6;necf6c2[1870]<=jcf1bb3;necf6c2[1852]<=jpf6dd6[0];necf6c2[1813]<=ou8d622;necf6c2[1799]<=uk10db8;necf6c2[1708]<=hq1bf36[0];necf6c2[1656]<=ri11ac4;necf6c2[1578]<=ng83d4e[0];necf6c2[1573]<=tudff4f;necf6c2[1551]<=ng86dc0;necf6c2[1493]<=en7f8df;necf6c2[1491]<=jrbfc6e;necf6c2[1417]<=mgb37fd;necf6c2[1396]<=ux26ff1[0];necf6c2[1378]<=xje6cdf[0];necf6c2[1368]<=vidf9b3[0];necf6c2[1353]<=jcc5f7a;necf6c2[1345]<=ui72605;necf6c2[1316]<=qg7de9b[0];necf6c2[1285]<=mg9814a[0];necf6c2[1265]<=ale2358;necf6c2[1198]<=bl7b137;necf6c2[1169]<=cz7a6c8;necf6c2[1163]<=ald9166;necf6c2[1117]<=kf2cd7f;necf6c2[1108]<=ba1ea72[0];necf6c2[1098]<=meffa7b;necf6c2[1054]<=cb36e02;necf6c2[1045]<=ym528b[0];necf6c2[1023]<=dmfe774;necf6c2[975]<=fc14694;necf6c2[965]<=shd6c1e[0];necf6c2[939]<=ldfc6fc;necf6c2[935]<=xwfe376;necf6c2[786]<=xl9bfe9;necf6c2[746]<=hdaff1b;necf6c2[745]<=bn37f8d;necf6c2[708]<=yz366ff;necf6c2[698]<=suc4dfe[0];necf6c2[689]<=fnfcd9b[0];necf6c2[676]<=tu58bef;necf6c2[672]<=ip4e4c0;necf6c2[658]<=zm2fbd3;necf6c2[642]<=hq93029;necf6c2[599]<=pf4f626[0];necf6c2[584]<=eaef4d9;necf6c2[581]<=vx9b22c;necf6c2[558]<=hb459af;necf6c2[522]<=jcc0a51[0];necf6c2[487]<=ux28d2;necf6c2[482]<=fpbad83[0];necf6c2[373]<=xy35fe3;necf6c2[349]<=rtd89bf;necf6c2[338]<=lf8b17d;necf6c2[336]<=lq58886;necf6c2[299]<=zxe9ec4[0];necf6c2[290]<=yxd3645;necf6c2[279]<=thc8b35;necf6c2[243]<=zkc051a;necf6c2[186]<=xw66bfc;necf6c2[169]<=gb5162f[0];necf6c2[168]<=wwc4432;necf6c2[149]<=wjfd3d8;necf6c2[121]<=twb80a3;necf6c2[84]<=th4a2c5[0];necf6c2[60]<=pub7014[0];necf6c2[42]<=mt29458[0];end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule