module s17;
 final begin
    $write("*-* All Finished *-*\n");
 end
endmodule