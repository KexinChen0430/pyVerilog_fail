module var_unnamed_block;
   initial begin
      integer var_in_unnamed;
   end
endmodule