module SCB_P4_v2_0_3 (
    interrupt,
    clock);
    output      interrupt;
    input       clock;
          wire  Net_904;
          wire  Net_898;
          wire  Net_933;
          wire  uncfg_rx_irq;
          wire  Net_824;
          wire  Net_823;
          wire  Net_767;
          wire  Net_754;
          wire  rx_irq;
          wire [3:0] ss;
          wire  Net_682;
          wire  Net_676;
          wire  Net_458;
          wire  Net_896;
          wire  Net_903;
          wire  Net_932;
          wire  Net_855;
          wire  Net_422;
          wire  Net_467;
          wire  SCBclock;
          wire  Net_751;
          wire  Net_928;
          wire  Net_927;
          wire  Net_459;
          wire  Net_747;
          wire  Net_746;
          wire  Net_452;
          wire  Net_379;
          wire  Net_654;
          wire  Net_416;
          wire  Net_891;
          wire  Net_387;
          wire  Net_653;
          wire  Net_739;
          wire  Net_916;
          wire  Net_660;
          wire  Net_915;
          wire  Net_252;
          wire  Net_899;
          wire  Net_652;
          wire  Net_474;
          wire  Net_909;
          wire  Net_547;
          wire  Net_245;
          wire  Net_663;
          wire  Net_847;
          wire  Net_656;
          wire  Net_703;
          wire  Net_687;
          wire  Net_581;
          wire  Net_580;
	cy_clock_v1_0
		#(.id("8c8734ef-3644-4eed-bc55-360072b94fff/81fcee8a-3b8b-4be1-9a5f-a5e2e619a938"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("62500000"),
		  .is_direct(0),
		  .is_digital(0))
		SCBCLK
		 (.clock_out(Net_847));
    ZeroTerminal ZeroTerminal_5 (
        .z(Net_459));
	wire [0:0] tmpOE__ss_s_net;
	wire [0:0] tmpIO_0__ss_s_net;
	wire [0:0] tmpINTERRUPT_0__ss_s_net;
	electrical [0:0] tmpSIOVREF__ss_s_net;
	cy_psoc3_pins_v1_10
		#(.id("8c8734ef-3644-4eed-bc55-360072b94fff/3446580a-3b9d-491c-8730-f7ea34ca86e3"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		ss_s
		 (.oe(tmpOE__ss_s_net),
		  .y({1'b0}),
		  .fb({Net_458}),
		  .io({tmpIO_0__ss_s_net[0:0]}),
		  .siovref(tmpSIOVREF__ss_s_net),
		  .interrupt({tmpINTERRUPT_0__ss_s_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__ss_s_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	// select_s_VM (cy_virtualmux_v1_0)
	assign Net_652 = Net_458;
    ZeroTerminal ZeroTerminal_4 (
        .z(Net_452));
    ZeroTerminal ZeroTerminal_3 (
        .z(Net_676));
    ZeroTerminal ZeroTerminal_2 (
        .z(Net_245));
    ZeroTerminal ZeroTerminal_1 (
        .z(Net_416));
	// rx_VM (cy_virtualmux_v1_0)
	assign Net_654 = Net_452;
	// rx_wake_VM (cy_virtualmux_v1_0)
	assign Net_682 = uncfg_rx_irq;
	// clock_VM (cy_virtualmux_v1_0)
	assign SCBclock = Net_847;
	// sclk_s_VM (cy_virtualmux_v1_0)
	assign Net_653 = Net_387;
	// mosi_s_VM (cy_virtualmux_v1_0)
	assign Net_909 = Net_252;
	// miso_m_VM (cy_virtualmux_v1_0)
	assign Net_663 = Net_245;
	wire [0:0] tmpOE__miso_s_net;
	wire [0:0] tmpFB_0__miso_s_net;
	wire [0:0] tmpIO_0__miso_s_net;
	wire [0:0] tmpINTERRUPT_0__miso_s_net;
	electrical [0:0] tmpSIOVREF__miso_s_net;
	cy_psoc3_pins_v1_10
		#(.id("8c8734ef-3644-4eed-bc55-360072b94fff/52f31aa9-2f0a-497d-9a1f-1424095e13e6"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("B"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		miso_s
		 (.oe(tmpOE__miso_s_net),
		  .y({Net_703}),
		  .fb({tmpFB_0__miso_s_net[0:0]}),
		  .io({tmpIO_0__miso_s_net[0:0]}),
		  .siovref(tmpSIOVREF__miso_s_net),
		  .interrupt({tmpINTERRUPT_0__miso_s_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__miso_s_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    ZeroTerminal ZeroTerminal_7 (
        .z(Net_754));
    assign Net_767 = Net_847 | Net_754;
	wire [0:0] tmpOE__sclk_s_net;
	wire [0:0] tmpIO_0__sclk_s_net;
	wire [0:0] tmpINTERRUPT_0__sclk_s_net;
	electrical [0:0] tmpSIOVREF__sclk_s_net;
	cy_psoc3_pins_v1_10
		#(.id("8c8734ef-3644-4eed-bc55-360072b94fff/4c15b41e-e284-4978-99e7-5aaee19bd0ce"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		sclk_s
		 (.oe(tmpOE__sclk_s_net),
		  .y({1'b0}),
		  .fb({Net_387}),
		  .io({tmpIO_0__sclk_s_net[0:0]}),
		  .siovref(tmpSIOVREF__sclk_s_net),
		  .interrupt({tmpINTERRUPT_0__sclk_s_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__sclk_s_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__mosi_s_net;
	wire [0:0] tmpIO_0__mosi_s_net;
	wire [0:0] tmpINTERRUPT_0__mosi_s_net;
	electrical [0:0] tmpSIOVREF__mosi_s_net;
	cy_psoc3_pins_v1_10
		#(.id("8c8734ef-3644-4eed-bc55-360072b94fff/5e2b647c-52cb-4f09-80bd-87ed9563ab24"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		mosi_s
		 (.oe(tmpOE__mosi_s_net),
		  .y({1'b0}),
		  .fb({Net_252}),
		  .io({tmpIO_0__mosi_s_net[0:0]}),
		  .siovref(tmpSIOVREF__mosi_s_net),
		  .interrupt({tmpINTERRUPT_0__mosi_s_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__mosi_s_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	// cts_VM (cy_virtualmux_v1_0)
	assign Net_739 = Net_747;
    cy_m0s8_scb_v2_0 SCB (
        .rx(Net_654),
        .miso_m(Net_663),
        .select_m(ss[3:0]),
        .sclk_m(Net_687),
        .mosi_s(Net_909),
        .select_s(Net_652),
        .sclk_s(Net_653),
        .mosi_m(Net_660),
        .scl(Net_580),
        .sda(Net_581),
        .tx(Net_656),
        .miso_s(Net_703),
        .interrupt(interrupt),
        .cts(Net_739),
        .rts(Net_751),
        .tx_req(Net_823),
        .rx_req(Net_824),
        .clock(SCBclock));
    defparam SCB.scb_mode = 1;
    ZeroTerminal ZeroTerminal_6 (
        .z(Net_747));
	// Device_VM1 (cy_virtualmux_v1_0)
	assign Net_547 = Net_896;
	// Device_VM5 (cy_virtualmux_v1_0)
	assign Net_891 = Net_932;
	// Device_VM2 (cy_virtualmux_v1_0)
	assign Net_474 = Net_903;
	// Device_VM3 (cy_virtualmux_v1_0)
	assign Net_899 = Net_915;
	// Device_VM4 (cy_virtualmux_v1_0)
	assign uncfg_rx_irq = Net_927;
endmodule