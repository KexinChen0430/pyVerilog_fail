module RESISTOR(1 2);
	parameter value=1;
	resistor #(.r(value)) r(1,2);
endmodule