module header
	// Internal signals
		// Generated Signal List
		// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances
	// wiring ...
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for i_avfb_tc_ctrl
		avfb_tc_ctrl i_avfb_tc_ctrl (
		);
		// End of Generated Instance Port Map for i_avfb_tc_ctrl
endmodule