module Test (
	     output wire out1 = 1'b1,
	     output integer out18 = 32'h18,
	     output var out1b = 1'b1,
	     output var logic out19 = 1'b1
	     );
endmodule