module IIR_Biquad_inj (clk,n_reset,sample_trig,X_in,filter_done,Y_out,p_desc86_p_O_FDE,p_desc87_p_O_FDE,p_desc88_p_O_FDE,p_desc89_p_O_FDE,p_desc90_p_O_FDE,p_desc91_p_O_FDE,p_desc92_p_O_FDE,p_desc93_p_O_FDE,p_desc94_p_O_FDE,p_desc95_p_O_FDE,p_desc96_p_O_FDE,p_desc97_p_O_FDE,p_desc98_p_O_FDE,p_desc99_p_O_FDE,p_desc100_p_O_FDE,p_desc101_p_O_FDE,p_desc102_p_O_FDE,p_desc103_p_O_FDE,p_desc104_p_O_FDE,p_desc105_p_O_FDE,p_desc106_p_O_FDE,p_desc107_p_O_FDE,p_desc108_p_O_FDE,p_desc109_p_O_FDE,p_desc110_p_O_FDE,p_desc111_p_O_FDE,p_desc112_p_O_FDE,p_desc113_p_O_FDE,p_desc114_p_O_FDE,p_desc115_p_O_FDE,p_desc116_p_O_FDE,p_desc117_p_O_FDE,p_desc118_p_O_FDE,p_desc119_p_O_FDE,p_desc120_p_O_FDE,p_desc121_p_O_FDE,p_desc162_p_O_FDE,p_desc163_p_O_FDE,p_desc164_p_O_FDE,p_desc165_p_O_FDE,p_desc166_p_O_FDE,p_desc167_p_O_FDE,p_desc168_p_O_FDE,p_desc169_p_O_FDE,p_desc170_p_O_FDE,p_desc171_p_O_FDE,p_desc172_p_O_FDE,p_desc173_p_O_FDE,p_desc174_p_O_FDE,p_desc175_p_O_FDE,p_desc176_p_O_FDE,p_desc177_p_O_FDE,p_desc178_p_O_FDE,p_desc179_p_O_FDE,p_desc198_p_O_FDE,p_desc199_p_O_FDE,p_desc200_p_O_FDE,p_desc201_p_O_FDE,p_desc202_p_O_FDE,p_desc203_p_O_FDE,p_desc204_p_O_FDE,p_desc205_p_O_FDE,p_desc206_p_O_FDE,p_desc207_p_O_FDE,p_desc208_p_O_FDE,p_desc209_p_O_FDE,p_desc210_p_O_FDE,p_desc211_p_O_FDE,p_desc212_p_O_FDE,p_desc213_p_O_FDE,p_desc214_p_O_FDE,p_desc215_p_O_FDE,p_desc216_p_O_FDE,p_desc217_p_O_FDE,p_desc218_p_O_FDE,p_desc219_p_O_FDE,p_desc220_p_O_FDE,p_desc221_p_O_FDE,p_desc222_p_O_FDE,p_desc223_p_O_FDE,p_desc224_p_O_FDE,p_desc225_p_O_FDE,p_desc226_p_O_FDE,p_desc227_p_O_FDE,p_desc228_p_O_FDE,p_desc229_p_O_FDE,p_desc230_p_O_FDE,p_desc231_p_O_FDE,p_desc232_p_O_FDE,p_desc233_p_O_FDE,p_desc234_p_O_FDE,p_desc235_p_O_FDE,p_desc236_p_O_FDE,p_desc237_p_O_FDE,p_desc238_p_O_FDE,p_desc239_p_O_FDE,p_desc240_p_O_FDE,p_desc241_p_O_FDE,p_desc242_p_O_FDE,p_desc243_p_O_FDE,p_desc244_p_O_FDE,p_desc245_p_O_FDE,p_desc246_p_O_FDE,p_desc247_p_O_FDE,p_desc248_p_O_FDE,p_desc249_p_O_FDE,p_desc250_p_O_FDE,p_desc251_p_O_FDE,p_desc252_p_O_FDE,p_desc253_p_O_FDE,p_desc254_p_O_FDE,p_desc255_p_O_FDE,p_desc256_p_O_FDE,p_desc257_p_O_FDE,p_desc258_p_O_FDE,p_desc259_p_O_FDE,p_desc260_p_O_FDE,p_desc261_p_O_FDE,p_desc262_p_O_FDE,p_desc263_p_O_FDE,p_desc264_p_O_FDE,p_desc334_p_O_FDC,p_desc335_p_O_FDC,p_desc336_p_O_FDC,p_desc337_p_O_FDC,p_state_reg_ret_5_Z_p_O_FDC,p_state_reg_ret_Z_p_O_FDP,p_state_reg_ret_1_Z_p_O_FDP,p_state_reg_ret_2_Z_p_O_FDP,p_state_reg_ret_4_Z_p_O_FDP,p_desc180_p_O_FDCE,p_desc181_p_O_FDCE,p_desc182_p_O_FDCE,p_desc183_p_O_FDCE,p_desc184_p_O_FDCE,p_desc185_p_O_FDCE,p_desc186_p_O_FDCE,p_desc187_p_O_FDCE,p_desc188_p_O_FDCE,p_desc189_p_O_FDCE,p_desc190_p_O_FDCE,p_desc191_p_O_FDCE,p_desc192_p_O_FDCE,p_desc193_p_O_FDCE,p_desc194_p_O_FDCE,p_desc195_p_O_FDCE,p_desc196_p_O_FDCE,p_desc197_p_O_FDCE,p_desc265_p_O_FDCE,p_desc266_p_O_FDCE,p_desc267_p_O_FDCE,p_desc268_p_O_FDCE,p_desc269_p_O_FDCE,p_desc270_p_O_FDCE,p_desc271_p_O_FDCE,p_desc272_p_O_FDCE,p_desc273_p_O_FDCE,p_desc274_p_O_FDCE,p_desc275_p_O_FDCE,p_desc276_p_O_FDCE,p_desc277_p_O_FDCE,p_desc278_p_O_FDCE,p_desc279_p_O_FDCE,p_desc280_p_O_FDCE,p_desc281_p_O_FDCE,p_desc282_p_O_FDCE,p_desc283_p_O_FDCE,p_desc284_p_O_FDCE,p_desc285_p_O_FDCE,p_desc286_p_O_FDCE,p_desc287_p_O_FDCE,p_desc288_p_O_FDCE,p_desc289_p_O_FDCE,p_desc290_p_O_FDCE,p_desc291_p_O_FDCE,p_desc292_p_O_FDCE,p_desc293_p_O_FDCE,p_desc294_p_O_FDCE,p_desc295_p_O_FDCE,p_desc296_p_O_FDCE,p_desc297_p_O_FDCE,p_desc298_p_O_FDCE,p_desc299_p_O_FDCE,p_desc300_p_O_FDCE,p_desc301_p_O_FDCE,p_desc302_p_O_FDCE,p_desc303_p_O_FDCE,p_desc304_p_O_FDCE,p_desc305_p_O_FDCE,p_desc306_p_O_FDCE,p_desc307_p_O_FDCE,p_desc308_p_O_FDCE,p_desc309_p_O_FDCE,p_desc310_p_O_FDCE,p_desc311_p_O_FDCE,p_desc312_p_O_FDCE,p_desc313_p_O_FDCE,p_desc314_p_O_FDCE,p_desc315_p_O_FDCE,p_desc316_p_O_FDCE,p_desc317_p_O_FDCE,p_desc318_p_O_FDCE,p_desc319_p_O_FDCE,p_desc320_p_O_FDCE,p_desc321_p_O_FDCE,p_desc322_p_O_FDCE,p_desc323_p_O_FDCE,p_desc324_p_O_FDCE,p_desc325_p_O_FDCE,p_desc326_p_O_FDCE,p_desc327_p_O_FDCE,p_desc328_p_O_FDCE,p_desc329_p_O_FDCE,p_desc330_p_O_FDCE,p_desc331_p_O_FDCE,p_desc332_p_O_FDCE,p_desc333_p_O_FDCE,p_desc338_p_O_FDCE,p_ZFF_Y1_0_rep1_Z_p_O_FDCE,p_desc339_p_O_FDCE,p_ZFF_Y1_15_rep1_Z_p_O_FDCE,p_desc340_p_O_FDCE,p_ZFF_X0_7_rep1_Z_p_O_FDCE,p_desc341_p_O_FDCE,p_desc342_p_O_FDCE,p_desc343_p_O_FDCE,p_desc344_p_O_FDCE,p_ZFF_Y1_16_rep1_Z_p_O_FDCE,p_desc345_p_O_FDCE,p_ZFF_X0_6_rep1_Z_p_O_FDCE,p_desc346_p_O_FDCE,p_desc347_p_O_FDCE,p_ZFF_Y1_2_rep1_Z_p_O_FDCE,p_desc348_p_O_FDCE,p_desc349_p_O_FDCE,p_ZFF_X0_10_rep1_Z_p_O_FDCE,p_desc350_p_O_FDCE,p_ZFF_X0_11_rep1_Z_p_O_FDCE,p_desc351_p_O_FDCE,p_ZFF_X0_12_rep1_Z_p_O_FDCE,p_desc352_p_O_FDCE,p_ZFF_X2_6_rep1_Z_p_O_FDCE,p_desc353_p_O_FDCE,p_ZFF_X0_4_rep1_Z_p_O_FDCE,p_desc354_p_O_FDCE,p_desc355_p_O_FDCE,p_desc356_p_O_FDCE,p_desc357_p_O_FDCE,p_ZFF_X2_10_rep1_Z_p_O_FDCE,p_desc358_p_O_FDCE,p_ZFF_X0_2_rep1_Z_p_O_FDCE,p_desc359_p_O_FDCE,p_ZFF_X0_1_rep1_Z_p_O_FDCE,p_desc360_p_O_FDCE,p_ZFF_Y1_1_rep1_Z_p_O_FDCE,p_desc361_p_O_FDCE,p_desc362_p_O_FDCE,p_desc363_p_O_FDCE,p_desc364_p_O_FDCE,p_ZFF_X2_2_rep1_Z_p_O_FDCE,p_desc365_p_O_FDCE,p_ZFF_X0_3_rep1_Z_p_O_FDCE,p_desc366_p_O_FDCE,p_desc367_p_O_FDCE,p_ZFF_X2_3_rep1_Z_p_O_FDCE,p_desc368_p_O_FDCE,p_ZFF_Y1_4_rep1_Z_p_O_FDCE,p_desc369_p_O_FDCE,p_desc370_p_O_FDCE,p_ZFF_Y1_3_rep1_Z_p_O_FDCE,p_desc371_p_O_FDCE,p_desc372_p_O_FDCE,p_desc373_p_O_FDCE,p_ZFF_Y1_5_rep1_Z_p_O_FDCE,p_desc374_p_O_FDCE,p_ZFF_X2_14_rep1_Z_p_O_FDCE,p_desc375_p_O_FDCE,p_ZFF_X0_14_rep1_Z_p_O_FDCE,p_desc376_p_O_FDCE,p_ZFF_X0_15_rep1_Z_p_O_FDCE,p_desc377_p_O_FDCE,p_ZFF_X2_15_rep1_Z_p_O_FDCE,p_desc378_p_O_FDCE,p_ZFF_Y1_6_rep1_Z_p_O_FDCE,p_desc379_p_O_FDCE,p_ZFF_Y1_13_rep1_Z_p_O_FDCE,p_desc380_p_O_FDCE,p_ZFF_Y1_7_rep1_Z_p_O_FDCE,p_desc381_p_O_FDCE,p_ZFF_Y1_14_rep1_Z_p_O_FDCE,p_desc382_p_O_FDCE,p_ZFF_X1_3_rep1_Z_p_O_FDCE,p_desc383_p_O_FDCE,p_ZFF_X1_0_rep1_Z_p_O_FDCE,p_desc384_p_O_FDCE,p_ZFF_Y1_9_rep1_Z_p_O_FDCE,p_desc385_p_O_FDCE,p_ZFF_X1_7_rep1_Z_p_O_FDCE,p_desc386_p_O_FDCE,p_ZFF_X1_4_rep1_Z_p_O_FDCE,p_desc387_p_O_FDCE,p_ZFF_X1_1_rep1_Z_p_O_FDCE,p_desc388_p_O_FDCE,p_ZFF_Y1_10_rep1_Z_p_O_FDCE,p_desc389_p_O_FDCE,p_ZFF_X1_8_rep1_Z_p_O_FDCE,p_desc390_p_O_FDCE,p_ZFF_X1_9_rep1_Z_p_O_FDCE,p_desc391_p_O_FDCE,p_ZFF_X1_11_rep1_Z_p_O_FDCE,p_desc392_p_O_FDCE,p_ZFF_X1_15_rep1_Z_p_O_FDCE,p_desc393_p_O_FDCE,p_ZFF_X1_2_rep1_Z_p_O_FDCE,p_desc394_p_O_FDCE,p_ZFF_Y1_12_rep1_Z_p_O_FDCE,p_desc395_p_O_FDCE,p_ZFF_X0_16_rep1_Z_p_O_FDCE,p_desc396_p_O_FDCE,p_desc397_p_O_FDCE,p_ZFF_Y1_17_rep1_Z_p_O_FDCE,p_desc398_p_O_FDCE,p_ZFF_X1_5_rep1_Z_p_O_FDCE,p_desc399_p_O_FDCE,p_ZFF_Y1_8_rep1_Z_p_O_FDCE,p_desc400_p_O_FDCE,p_desc401_p_O_FDCE,p_desc402_p_O_FDCE,p_ZFF_X1_6_rep1_Z_p_O_FDCE,p_desc403_p_O_FDCE,p_ZFF_X1_12_rep1_Z_p_O_FDCE,p_desc404_p_O_FDCE,p_ZFF_X1_10_rep1_Z_p_O_FDCE,p_desc405_p_O_FDCE,p_ZFF_X1_13_rep1_Z_p_O_FDCE,p_desc406_p_O_FDCE,p_ZFF_Y1_11_rep1_Z_p_O_FDCE,p_desc407_p_O_FDCE,p_ZFF_Y2_8_rep1_Z_p_O_FDCE,p_desc408_p_O_FDCE,p_desc409_p_O_FDCE,p_ZFF_Y2_6_rep1_Z_p_O_FDCE,p_desc410_p_O_FDCE,p_ZFF_Y2_7_rep1_Z_p_O_FDCE,p_desc411_p_O_FDCE,p_ZFF_Y2_14_rep1_Z_p_O_FDCE);
input clk ;
input n_reset ;
input sample_trig ;
input [17:0] X_in ;
output filter_done ;
output [17:0] Y_out ;
wire clk ;
wire n_reset ;
wire sample_trig ;
wire filter_done ;
wire [2:0] q_reg ;
wire [17:0] pgZFF_Y1 ;
wire [17:0] pgZFF_Y2 ;
wire [16:0] ZFF_X0 ;
wire [17:0] ZFF_Y2 ;
wire [42:8] un9_10 ;
wire [17:3] ZFF_Y1 ;
wire [46:22] un9_11 ;
wire [16:0] ZFF_X1 ;
wire [16:0] ZFF_X2 ;
wire state_reg ;
wire state_next ;
wire [46:30] pgZFF_X0_quad ;
wire [47:30] pgZFF_X1_quad ;
wire [46:30] pgZFF_X2_quad ;
wire [47:30] pgZFF_Y1_quad ;
wire [47:30] pgZFF_Y2_quad ;
wire [2:0] q_next ;
wire [16:0] pgZFF_X0 ;
wire [16:0] pgZFF_X2 ;
wire [17:0] pgZFF_X1 ;
wire [17:0] Y_out_double_2 ;
wire [17:0] Y_out_double ;
wire [2:0] q_reg_i_1 ;
wire [42:15] un6_0_9 ;
wire [39:10] un6_0_8 ;
wire [28:5] un6_0_6 ;
wire [45:18] un7_0_10 ;
wire [38:9] un7_0_8 ;
wire [33:3] un7_0_6 ;
wire [42:15] un8_0_9 ;
wire [39:10] un8_0_8 ;
wire [28:5] un8_0_6 ;
wire [36:6] un10_6 ;
wire [46:6] un9_8 ;
wire [47:2] un9_6 ;
wire [17:2] Y_out_double_2_7 ;
wire [17:0] Y_out_double_2_4 ;
wire [47:15] un10_8 ;
wire [17:0] Y_out_double_2_6 ;
wire [2:0] q_next_i ;
wire [1:1] pgZFF_X0_i ;
wire [17:17] un7_0_10_i_i ;
wire [47:44] un10_8_i ;
wire [6:6] un10_6_i ;
wire [23:23] un9_11_i ;
wire pgZFF_Y1_i ;
wire [8:8] un9_10_fast ;
wire [17:3] ZFF_Y1_fast ;
wire [16:0] ZFF_X0_fast ;
wire [16:0] ZFF_X2_fast ;
wire [7:6] un9_8_fast ;
wire [26:22] un9_11_fast ;
wire [16:0] ZFF_X1_fast ;
wire [17:6] ZFF_Y2_fast ;
wire [28:28] un6_0_6_0 ;
wire [28:28] un6_0_6_1 ;
wire [47:47] un9_6_0 ;
wire [47:47] un9_6_1 ;
wire [46:46] un9_8_1 ;
wire [42:42] un9_10_0 ;
wire [42:42] un9_10_1 ;
wire [36:36] un10_6_0 ;
wire [36:36] un10_6_1 ;
wire [28:28] un8_0_6_0 ;
wire [28:28] un8_0_6_1 ;
wire [33:33] un7_0_6_0 ;
wire [33:33] un7_0_6_1 ;
wire [38:38] un7_0_8_0 ;
wire [38:38] un7_0_8_1 ;
wire [39:39] un6_0_8_1 ;
wire [39:39] un8_0_8_1 ;
wire [42:42] un6_0_9_0 ;
wire [42:42] un6_0_9_1 ;
wire [42:42] un8_0_9_0 ;
wire [42:42] un8_0_9_1 ;
wire [46:46] un9_11_0 ;
wire [46:46] un9_11_1 ;
wire VCC ;
wire GND ;
wire state_reg_ret_4 ;
wire un7_0_0_s_29 ;
wire un7_0_0_s_30 ;
wire un7_0_0_s_31 ;
wire un7_0_0_s_32 ;
wire un7_0_0_s_33 ;
wire un7_0_0_s_34 ;
wire un7_0_0_s_35 ;
wire un7_0_0_s_36 ;
wire un7_0_0_s_37 ;
wire un7_0_0_s_38 ;
wire un7_0_0_s_39 ;
wire un7_0_0_s_40 ;
wire un7_0_0_s_41 ;
wire un7_0_0_s_42 ;
wire un7_0_0_s_43 ;
wire un7_0_0_s_44 ;
wire un7_0_0_s_45 ;
wire state_reg_ret_5_cb ;
wire sum_stg_a ;
wire trunc_out ;
wire trunc_prods ;
wire un7_q_reg_reti ;
wire un1_q_reg_2_reti ;
wire N_40 ;
wire N_371 ;
wire N_372 ;
wire N_373 ;
wire N_374 ;
wire un1_q_reg_2_c ;
wire un10_8_o5_11 ;
wire un10_8_o5_12 ;
wire un10_8_o5_13 ;
wire un10_8_o5_14 ;
wire un10_8_o5_15 ;
wire un10_8_o5_16 ;
wire un10_8_o5_17 ;
wire un10_8_o5_18 ;
wire un10_8_o5_19 ;
wire un10_8_o5_20 ;
wire un10_8_o5_21 ;
wire un10_8_o5_22 ;
wire un10_8_o5_23 ;
wire un8_0_8_cry_3_RNO ;
wire un8_0_8_cry_4_RNO ;
wire un8_0_8_o5_4 ;
wire un8_0_8_cry_6_RNO ;
wire un8_0_8_cry_7_RNO ;
wire un8_0_8_cry_8_RNO ;
wire un8_0_8_cry_9_RNO ;
wire un8_0_8_cry_10_RNO ;
wire un8_0_8_o5_10 ;
wire un8_0_8_o5_11 ;
wire un8_0_8_cry_13_RNO ;
wire un8_0_8_cry_14_RNO ;
wire un8_0_8_cry_16_RNO ;
wire un8_0_8_cry_18_RNO ;
wire un8_0_8_cry_20_RNO ;
wire un6_0_8_cry_3_RNO ;
wire un6_0_8_cry_4_RNO ;
wire un6_0_8_o5_4 ;
wire un6_0_8_cry_6_RNO ;
wire un6_0_8_cry_7_RNO ;
wire un6_0_8_cry_8_RNO ;
wire un6_0_8_cry_9_RNO ;
wire un6_0_8_cry_10_RNO ;
wire un6_0_8_o5_10 ;
wire un6_0_8_o5_11 ;
wire un6_0_8_cry_13_RNO ;
wire un6_0_8_cry_14_RNO ;
wire un6_0_8_cry_16_RNO ;
wire un6_0_8_cry_18_RNO ;
wire un6_0_8_cry_20_RNO ;
wire un7_0_8_cry_6_RNO ;
wire un7_0_8_cry_7_RNO ;
wire un7_0_8_cry_8_RNO ;
wire un7_0_8_cry_9_RNO ;
wire un7_0_8_cry_10_RNO ;
wire un7_0_8_cry_11_RNO ;
wire un7_0_8_cry_12_RNO ;
wire un7_0_8_cry_13_RNO ;
wire un7_0_8_cry_14_RNO ;
wire un7_0_8_cry_15_RNO ;
wire un7_0_8_cry_16_RNO ;
wire un7_0_8_cry_17_RNO ;
wire un7_0_8_cry_18_RNO ;
wire un7_0_8_cry_19_RNO ;
wire un7_0_6_cry_5_RNO ;
wire un7_0_6_cry_10_RNO ;
wire un7_0_6_cry_11_RNO ;
wire un7_0_6_cry_12_RNO ;
wire un7_0_6_cry_13_RNO ;
wire un7_0_6_cry_14_RNO ;
wire un7_0_6_cry_15_RNO ;
wire un7_0_6_o5_15 ;
wire un7_0_6_o5_16 ;
wire un7_0_6_o5_17 ;
wire un7_0_6_o5_18 ;
wire un7_0_6_o5_19 ;
wire un7_0_6_o5_20 ;
wire un7_0_6_cry_22_RNO ;
wire un7_0_0_axb_10_lut6_2_O5 ;
wire un7_0_0_o5_11 ;
wire un7_0_0_o5_12 ;
wire un7_0_0_o5_13 ;
wire un7_0_0_o5_14 ;
wire un7_0_0_o5_15 ;
wire un7_0_0_o5_16 ;
wire un7_0_0_o5_17 ;
wire un7_0_0_o5_18 ;
wire un7_0_0_o5_19 ;
wire un7_0_0_o5_20 ;
wire un7_0_0_o5_21 ;
wire un7_0_0_o5_22 ;
wire un7_0_0_o5_23 ;
wire un7_0_0_o5_24 ;
wire un7_0_0_o5_25 ;
wire un7_0_0_o5_26 ;
wire un7_0_0_o5_27 ;
wire un7_0_0_o5_28 ;
wire un7_0_0_o5_29 ;
wire un7_0_0_o5_30 ;
wire un7_0_0_o5_31 ;
wire un7_0_0_o5_32 ;
wire un7_0_0_cry_34_RNO ;
wire un7_0_0_cry_39_RNO ;
wire un8_0_6_1_scalar ;
wire un8_0_6_cry_5_RNO ;
wire un8_0_6_cry_6_RNO ;
wire un8_0_6_cry_7_RNO ;
wire un8_0_6_cry_8_RNO ;
wire un8_0_6_cry_9_RNO ;
wire un8_0_6_cry_10_RNO ;
wire un8_0_6_cry_11_RNO ;
wire un8_0_6_cry_12_RNO ;
wire un8_0_6_cry_13_RNO ;
wire un8_0_6_cry_14_RNO ;
wire un8_0_6_cry_15_RNO ;
wire un8_0_6_cry_16_RNO ;
wire un8_0_6_cry_17_RNO ;
wire un8_0_6_cry_18_RNO ;
wire un8_0_6_cry_19_RNO ;
wire un8_0_0_axb_11_lut6_2_O5 ;
wire un8_0_0_o5_12 ;
wire un8_0_0_o5_13 ;
wire un8_0_0_o5_14 ;
wire un8_0_0_o5_15 ;
wire un8_0_0_o5_16 ;
wire un8_0_0_o5_17 ;
wire un8_0_0_o5_18 ;
wire un8_0_0_o5_19 ;
wire un8_0_0_o5_20 ;
wire un8_0_0_o5_21 ;
wire un8_0_0_o5_22 ;
wire un8_0_0_o5_23 ;
wire un8_0_0_o5_24 ;
wire un8_0_0_o5_25 ;
wire un8_0_0_o5_26 ;
wire un8_0_0_o5_27 ;
wire un8_0_0_cry_29_RNO ;
wire un8_0_8_s_26_RNIUCD71_O5 ;
wire un8_0_0_o5_37 ;
wire un8_0_0_o5_41 ;
wire un10_6_cry_0_RNO ;
wire un10_6_cry_4_RNO ;
wire un10_6_cry_5_RNO ;
wire un10_6_cry_6_RNO ;
wire un10_6_cry_7_RNO ;
wire un10_6_cry_8_RNO ;
wire un10_6_cry_9_RNO ;
wire un10_6_cry_10_RNO ;
wire un10_6_cry_11_RNO ;
wire un10_6_cry_12_RNO ;
wire un10_6_cry_13_RNO ;
wire un10_6_cry_14_RNO ;
wire un10_6_cry_15_RNO ;
wire un10_6_cry_16_RNO ;
wire un10_6_cry_17_RNO ;
wire un10_6_cry_18_RNO ;
wire un10_6_cry_19_RNO ;
wire un10_6_cry_20_RNO ;
wire un10_10 ;
wire un10_19 ;
wire un10_29 ;
wire un10_axb_11_lut6_2_O5 ;
wire un10_o5_12 ;
wire un10_o5_13 ;
wire un10_o5_14 ;
wire un10_o5_15 ;
wire un10_o5_16 ;
wire un10_o5_17 ;
wire un10_o5_18 ;
wire un10_o5_19 ;
wire un10_o5_20 ;
wire un10_o5_21 ;
wire un10_o5_22 ;
wire un10_o5_23 ;
wire un10_o5_24 ;
wire un10_o5_25 ;
wire un10_o5_26 ;
wire un10_o5_27 ;
wire un10_cry_29_RNO ;
wire un10_cry_31_RNO ;
wire un9_10_cry_3_RNO ;
wire un9_10_cry_6_RNO ;
wire un9_10_cry_7_RNO ;
wire un9_10_cry_9_RNO ;
wire un9_10_cry_10_RNO ;
wire un9_10_cry_11_RNO ;
wire un9_10_cry_12_RNO ;
wire un9_10_cry_13_RNO ;
wire un9_10_cry_14_RNO ;
wire un9_10_cry_15_RNO ;
wire un9_10_cry_16_RNO ;
wire un9_10_cry_17_RNO ;
wire un9_10_cry_18_RNO ;
wire un9_10_cry_19_RNO ;
wire un9_10_cry_20_RNO ;
wire un9_10_cry_21_RNO ;
wire un9_10_cry_22_RNO ;
wire un9_10_cry_23_RNO ;
wire un9_10_cry_24_RNO ;
wire un9_8_cry_7_RNO ;
wire un9_8_cry_8_RNO ;
wire un9_8_cry_9_RNO ;
wire un9_8_cry_10_RNO ;
wire un9_8_cry_11_RNO ;
wire un9_8_cry_12_RNO ;
wire un9_8_cry_13_RNO ;
wire un9_8_o5_13 ;
wire un9_8_o5_14 ;
wire un9_8_o5_15 ;
wire un9_8_cry_17_RNO ;
wire un9_8_o5_17 ;
wire un9_8_o5_18 ;
wire un9_8_o5_19 ;
wire un9_8_cry_21_RNO ;
wire un9_6_0_cry_6_RNO ;
wire un9_6_0_cry_7_RNO ;
wire un9_6_0_cry_8_RNO ;
wire un9_6_0_cry_11_RNO ;
wire un9_6_0_cry_12_RNO ;
wire un9_6_0_cry_13_RNO ;
wire un9_6_0_cry_14_RNO ;
wire un9_6_0_cry_15_RNO ;
wire un9_6_0_cry_16_RNO ;
wire un9_6_0_cry_17_RNO ;
wire un9_6_0_cry_18_RNO ;
wire un9_6_0_cry_19_RNO ;
wire un9_6_0_cry_20_RNO ;
wire un9_6_78 ;
wire un9_6_0_cry_22_RNO ;
wire un9_6_0_cry_23_RNO ;
wire un9_6_0_cry_24_RNO ;
wire un9_6_0_cry_25_RNO ;
wire un9_6_0_cry_26_RNO ;
wire un9_6_0_cry_27_RNO ;
wire un9_6_0_cry_28_RNO ;
wire un9_6_0_cry_29_RNO ;
wire un9_6_0_cry_31_RNO ;
wire un9_o5_7 ;
wire un9_o5_8 ;
wire un9_o5_9 ;
wire un9_o5_10 ;
wire un9_o5_11 ;
wire un9_o5_12 ;
wire un9_o5_13 ;
wire un9_o5_14 ;
wire un9_o5_15 ;
wire un9_o5_16 ;
wire un9_o5_17 ;
wire un9_o5_18 ;
wire un9_o5_19 ;
wire un9_o5_20 ;
wire un9_o5_21 ;
wire un9_o5_22 ;
wire un9_o5_23 ;
wire un9_o5_24 ;
wire un9_o5_25 ;
wire un9_o5_26 ;
wire un9_o5_27 ;
wire un9_o5_28 ;
wire un9_o5_29 ;
wire un9_o5_30 ;
wire un9_o5_31 ;
wire un9_o5_32 ;
wire un9_o5_33 ;
wire un9_o5_34 ;
wire un9_o5_35 ;
wire un9_o5_36 ;
wire un9_o5_37 ;
wire un9_o5_38 ;
wire un9_o5_39 ;
wire un9_cry_41_RNO ;
wire Y_out_double_2_6_0_o5_1 ;
wire Y_out_double_2_6_0_o5_2 ;
wire Y_out_double_2_6_0_o5_3 ;
wire Y_out_double_2_6_0_o5_4 ;
wire Y_out_double_2_6_0_o5_5 ;
wire Y_out_double_2_6_0_o5_6 ;
wire Y_out_double_2_6_0_o5_7 ;
wire Y_out_double_2_6_0_o5_8 ;
wire Y_out_double_2_6_0_o5_9 ;
wire Y_out_double_2_6_0_o5_10 ;
wire Y_out_double_2_6_0_o5_11 ;
wire Y_out_double_2_6_0_o5_12 ;
wire Y_out_double_2_6_0_o5_13 ;
wire Y_out_double_2_6_0_o5_14 ;
wire Y_out_double_2_6_0_o5_15 ;
wire un6_0_6_1_scalar ;
wire un6_0_6_cry_5_RNO ;
wire un6_0_6_cry_6_RNO ;
wire un6_0_6_cry_7_RNO ;
wire un6_0_6_cry_8_RNO ;
wire un6_0_6_cry_9_RNO ;
wire un6_0_6_cry_10_RNO ;
wire un6_0_6_cry_11_RNO ;
wire un6_0_6_cry_12_RNO ;
wire un6_0_6_cry_13_RNO ;
wire un6_0_6_cry_14_RNO ;
wire un6_0_6_cry_15_RNO ;
wire un6_0_6_cry_16_RNO ;
wire un6_0_6_cry_17_RNO ;
wire un6_0_6_cry_18_RNO ;
wire un6_0_6_cry_19_RNO ;
wire un6_0_0_axb_11_lut6_2_O5 ;
wire un6_0_0_o5_12 ;
wire un6_0_0_o5_13 ;
wire un6_0_0_o5_14 ;
wire un6_0_0_o5_15 ;
wire un6_0_0_o5_16 ;
wire un6_0_0_o5_17 ;
wire un6_0_0_o5_18 ;
wire un6_0_0_o5_19 ;
wire un6_0_0_o5_20 ;
wire un6_0_0_o5_21 ;
wire un6_0_0_o5_22 ;
wire un6_0_0_o5_23 ;
wire un6_0_0_o5_24 ;
wire un6_0_0_o5_25 ;
wire un6_0_0_o5_26 ;
wire un6_0_0_o5_27 ;
wire un6_0_0_cry_29_RNO ;
wire un6_0_9_s_21_RNIM4BU_O5 ;
wire un6_0_0_o5_37 ;
wire un6_0_0_o5_41 ;
wire un7_0_10_cry_0_RNO ;
wire un7_0_10_cry_14_RNO ;
wire un7_0_10_o5_14 ;
wire un7_0_10_o5_15 ;
wire un7_0_10_o5_16 ;
wire un7_0_10_14 ;
wire un7_0_10_o5_17 ;
wire un7_0_10_o5_18 ;
wire un7_0_10_o5_19 ;
wire un7_0_10_o5_20 ;
wire un7_0_10_o5_21 ;
wire un10_8_ac0_5 ;
wire un9_ac0_105 ;
wire un7_0_10_cry_0 ;
wire un7_0_10_cry_1_RNO ;
wire un7_0_10_axb_1 ;
wire un7_0_10_cry_1 ;
wire un7_0_10_axb_2 ;
wire un7_0_10_cry_2 ;
wire un7_0_10_axb_3 ;
wire un7_0_10_cry_3 ;
wire un7_0_10_axb_4 ;
wire un7_0_10_cry_4 ;
wire un7_0_10_axb_5 ;
wire un7_0_10_cry_5 ;
wire un7_0_10_axb_6 ;
wire un7_0_10_cry_6 ;
wire un7_0_10_axb_7 ;
wire un7_0_10_cry_7 ;
wire un7_0_10_axb_8 ;
wire un7_0_10_cry_8 ;
wire un7_0_10_axb_9 ;
wire un7_0_10_cry_9 ;
wire un7_0_10_axb_10 ;
wire un7_0_10_cry_10 ;
wire un7_0_10_axb_11 ;
wire un7_0_10_cry_11 ;
wire un7_0_10_cry_12_RNO ;
wire un7_0_10_axb_12 ;
wire un7_0_10_cry_12 ;
wire un7_0_10_cry_13_RNO ;
wire un7_0_10_axb_13 ;
wire un7_0_10_cry_13 ;
wire un7_0_10_axb_14 ;
wire un7_0_10_cry_14 ;
wire un7_0_10_axb_15 ;
wire un7_0_10_cry_15 ;
wire un7_0_10_axb_16 ;
wire un7_0_10_cry_16 ;
wire un7_0_10_axb_17 ;
wire un7_0_10_cry_17 ;
wire un7_0_10_axb_18 ;
wire un7_0_10_cry_18 ;
wire un7_0_10_axb_19 ;
wire un7_0_10_cry_19 ;
wire un7_0_10_axb_20 ;
wire un7_0_10_cry_20 ;
wire un7_0_10_axb_21 ;
wire un7_0_10_cry_21 ;
wire un7_0_10_axb_22 ;
wire un7_0_10_cry_22 ;
wire un7_0_10_axb_23 ;
wire un7_0_10_cry_23 ;
wire un7_0_10_cry_24 ;
wire un7_0_10_cry_25 ;
wire un7_0_10_axb_26 ;
wire un7_0_10_cry_26 ;
wire un6_0_0_s_28 ;
wire un6_0_0_s_29 ;
wire un6_0_0_s_30 ;
wire un6_0_0_s_31 ;
wire un6_0_0_s_32 ;
wire un6_0_0_s_33 ;
wire un6_0_0_s_34 ;
wire un6_0_0_s_35 ;
wire un6_0_0_s_36 ;
wire un6_0_0_s_37 ;
wire un6_0_0_s_38 ;
wire un6_0_0_s_39 ;
wire un6_0_0_s_40 ;
wire un6_0_0_s_41 ;
wire un6_0_0_s_42 ;
wire un6_0_0_s_43 ;
wire un6_0_0_cry_0 ;
wire un6_0_0_cry_1 ;
wire un6_0_0_cry_2 ;
wire un6_0_0_cry_3 ;
wire un6_0_0_cry_4 ;
wire un6_0_0_cry_5 ;
wire un6_0_0_cry_6 ;
wire un6_0_0_axb_7 ;
wire un6_0_0_cry_7 ;
wire un6_0_0_axb_8 ;
wire un6_0_0_cry_8 ;
wire un6_0_0_axb_9 ;
wire un6_0_0_cry_9 ;
wire un6_0_0_axb_10 ;
wire un6_0_0_cry_10 ;
wire un6_0_0_axb_11 ;
wire un6_0_0_cry_11 ;
wire un6_0_0_axb_12 ;
wire un6_0_0_cry_12 ;
wire un6_0_0_axb_13 ;
wire un6_0_0_cry_13 ;
wire un6_0_0_axb_14 ;
wire un6_0_0_cry_14 ;
wire un6_0_0_axb_15 ;
wire un6_0_0_cry_15 ;
wire un6_0_0_axb_16 ;
wire un6_0_0_cry_16 ;
wire un6_0_0_axb_17 ;
wire un6_0_0_cry_17 ;
wire un6_0_0_axb_18 ;
wire un6_0_0_cry_18 ;
wire un6_0_0_axb_19 ;
wire un6_0_0_cry_19 ;
wire un6_0_0_axb_20 ;
wire un6_0_0_cry_20 ;
wire un6_0_0_axb_21 ;
wire un6_0_0_cry_21 ;
wire un6_0_0_axb_22 ;
wire un6_0_0_cry_22 ;
wire un6_0_0_axb_23 ;
wire un6_0_0_cry_23 ;
wire un6_0_0_axb_24 ;
wire un6_0_0_cry_24 ;
wire un6_0_0_axb_25 ;
wire un6_0_0_cry_25 ;
wire un6_0_0_axb_26 ;
wire un6_0_0_cry_26 ;
wire un6_0_0_axb_27 ;
wire un6_0_0_cry_27 ;
wire un6_0_0_axb_28 ;
wire un6_0_0_cry_28 ;
wire un6_0_0_axb_29 ;
wire un6_0_0_cry_29 ;
wire un6_0_0_cry_30_RNO ;
wire un6_0_0_axb_30 ;
wire un6_0_0_cry_30 ;
wire un6_0_0_cry_31_RNO ;
wire un6_0_0_axb_31 ;
wire un6_0_0_cry_31 ;
wire un6_0_0_cry_32_RNO ;
wire un6_0_0_axb_32 ;
wire un6_0_0_cry_32 ;
wire un6_0_0_cry_33_RNO ;
wire un6_0_0_axb_33 ;
wire un6_0_0_cry_33 ;
wire un6_0_0_cry_34_RNO ;
wire un6_0_0_axb_34 ;
wire un6_0_0_cry_34 ;
wire un6_0_0_cry_35_RNO ;
wire un6_0_0_axb_35 ;
wire un6_0_0_cry_35 ;
wire un6_0_0_cry_36_RNO ;
wire un6_0_0_axb_36 ;
wire un6_0_0_cry_36 ;
wire un6_0_0_axb_37 ;
wire un6_0_0_cry_37 ;
wire un6_0_0_axb_38 ;
wire un6_0_0_cry_38 ;
wire un6_0_0_axb_39 ;
wire un6_0_0_cry_39 ;
wire un6_0_0_cry_40 ;
wire un6_0_0_axb_41 ;
wire un6_0_0_cry_41 ;
wire un6_0_0_axb_42 ;
wire un6_0_0_cry_42 ;
wire un6_0_0_axb_43 ;
wire un6_0_6_cry_0 ;
wire un6_0_6_axb_1 ;
wire un6_0_6_cry_1 ;
wire un6_0_6_axb_2 ;
wire un6_0_6_cry_2 ;
wire un6_0_6_axb_3 ;
wire un6_0_6_cry_3 ;
wire un6_0_6_cry_4_RNO ;
wire un6_0_6_axb_4 ;
wire un6_0_6_cry_4 ;
wire un6_0_6_axb_5 ;
wire un6_0_6_cry_5 ;
wire un6_0_6_axb_6 ;
wire un6_0_6_cry_6 ;
wire un6_0_6_axb_7 ;
wire un6_0_6_cry_7 ;
wire un6_0_6_axb_8 ;
wire un6_0_6_cry_8 ;
wire un6_0_6_axb_9 ;
wire un6_0_6_cry_9 ;
wire un6_0_6_axb_10 ;
wire un6_0_6_cry_10 ;
wire un6_0_6_axb_11 ;
wire un6_0_6_cry_11 ;
wire un6_0_6_axb_12 ;
wire un6_0_6_cry_12 ;
wire un6_0_6_axb_13 ;
wire un6_0_6_cry_13 ;
wire un6_0_6_axb_14 ;
wire un6_0_6_cry_14 ;
wire un6_0_6_axb_15 ;
wire un6_0_6_cry_15 ;
wire un6_0_6_axb_16 ;
wire un6_0_6_cry_16 ;
wire un6_0_6_axb_17 ;
wire un6_0_6_cry_17 ;
wire un6_0_6_axb_18 ;
wire un6_0_6_cry_18 ;
wire un6_0_6_axb_19 ;
wire un6_0_6_cry_19 ;
wire un6_0_6_cry_20_RNO ;
wire un6_0_6_axb_20 ;
wire un6_0_6_cry_20 ;
wire un6_0_6_43 ;
wire un6_0_6_axb_21 ;
wire un6_0_6_cry_21 ;
wire un6_0_6_axb_22 ;
wire Y_out_double_2_6_0_axb_0 ;
wire Y_out_double_2_6_0_cry_0 ;
wire Y_out_double_2_6_0_axb_1 ;
wire Y_out_double_2_6_0_cry_1 ;
wire Y_out_double_2_6_0_axb_2 ;
wire Y_out_double_2_6_0_cry_2 ;
wire Y_out_double_2_6_0_axb_3 ;
wire Y_out_double_2_6_0_cry_3 ;
wire Y_out_double_2_6_0_axb_4 ;
wire Y_out_double_2_6_0_cry_4 ;
wire Y_out_double_2_6_0_axb_5 ;
wire Y_out_double_2_6_0_cry_5 ;
wire Y_out_double_2_6_0_axb_6 ;
wire Y_out_double_2_6_0_cry_6 ;
wire Y_out_double_2_6_0_axb_7 ;
wire Y_out_double_2_6_0_cry_7 ;
wire Y_out_double_2_6_0_axb_8 ;
wire Y_out_double_2_6_0_cry_8 ;
wire Y_out_double_2_6_0_axb_9 ;
wire Y_out_double_2_6_0_cry_9 ;
wire Y_out_double_2_6_0_axb_10 ;
wire Y_out_double_2_6_0_cry_10 ;
wire Y_out_double_2_6_0_axb_11 ;
wire Y_out_double_2_6_0_cry_11 ;
wire Y_out_double_2_6_0_axb_12 ;
wire Y_out_double_2_6_0_cry_12 ;
wire Y_out_double_2_6_0_axb_13 ;
wire Y_out_double_2_6_0_cry_13 ;
wire Y_out_double_2_6_0_axb_14 ;
wire Y_out_double_2_6_0_cry_14 ;
wire Y_out_double_2_6_0_axb_15 ;
wire Y_out_double_2_6_0_cry_15 ;
wire Y_out_double_2_6_0_axb_16 ;
wire Y_out_double_2_6_0_cry_16 ;
wire Y_out_double_2_6_0_axb_17 ;
wire un9_s_28 ;
wire un9_s_29 ;
wire un9_s_30 ;
wire un9_s_31 ;
wire un9_s_32 ;
wire un9_s_33 ;
wire un9_s_34 ;
wire un9_s_35 ;
wire un9_s_36 ;
wire un9_s_37 ;
wire un9_s_38 ;
wire un9_s_39 ;
wire un9_s_40 ;
wire un9_s_41 ;
wire un9_s_42 ;
wire un9_s_43 ;
wire un9_s_44 ;
wire un9_s_45 ;
wire un9_cry_0 ;
wire un9_axb_1 ;
wire un9_cry_1 ;
wire un9_axb_2 ;
wire un9_cry_2 ;
wire un9_axb_3 ;
wire un9_cry_3 ;
wire un9_axb_4 ;
wire un9_cry_4 ;
wire un9_axb_5 ;
wire un9_cry_5 ;
wire un9_axb_6 ;
wire un9_cry_6 ;
wire un9_cry_7_RNO ;
wire un9_axb_7 ;
wire un9_cry_7 ;
wire un9_axb_8 ;
wire un9_cry_8 ;
wire un9_axb_9 ;
wire un9_cry_9 ;
wire un9_axb_10 ;
wire un9_cry_10 ;
wire un9_axb_11 ;
wire un9_cry_11 ;
wire un9_axb_12 ;
wire un9_cry_12 ;
wire un9_axb_13 ;
wire un9_cry_13 ;
wire un9_axb_14 ;
wire un9_cry_14 ;
wire un9_axb_15 ;
wire un9_cry_15 ;
wire un9_axb_16 ;
wire un9_cry_16 ;
wire un9_axb_17 ;
wire un9_cry_17 ;
wire un9_axb_18 ;
wire un9_cry_18 ;
wire un9_axb_19 ;
wire un9_cry_19 ;
wire un9_axb_20 ;
wire un9_cry_20 ;
wire un9_axb_21 ;
wire un9_cry_21 ;
wire un9_axb_22 ;
wire un9_cry_22 ;
wire un9_axb_23 ;
wire un9_cry_23 ;
wire un9_axb_24 ;
wire un9_cry_24 ;
wire un9_axb_25 ;
wire un9_cry_25 ;
wire un9_axb_26 ;
wire un9_cry_26 ;
wire un9_axb_27 ;
wire un9_cry_27 ;
wire un9_axb_28 ;
wire un9_cry_28 ;
wire un9_axb_29 ;
wire un9_cry_29 ;
wire un9_axb_30 ;
wire un9_cry_30 ;
wire un9_axb_31 ;
wire un9_cry_31 ;
wire un9_axb_32 ;
wire un9_cry_32 ;
wire un9_axb_33 ;
wire un9_cry_33 ;
wire un9_axb_34 ;
wire un9_cry_34 ;
wire un9_axb_35 ;
wire un9_cry_35 ;
wire un9_axb_36 ;
wire un9_cry_36 ;
wire un9_axb_37 ;
wire un9_cry_37 ;
wire un9_axb_38 ;
wire un9_cry_38 ;
wire un9_axb_39 ;
wire un9_cry_39 ;
wire un9_axb_40 ;
wire un9_cry_40 ;
wire un9_axb_41 ;
wire un9_cry_41 ;
wire un9_cry_42_RNO ;
wire un9_axb_42 ;
wire un9_cry_42 ;
wire un9_cry_43_RNO ;
wire un9_axb_43 ;
wire un9_cry_43 ;
wire un9_cry_44_RNO ;
wire un9_axb_44 ;
wire un9_cry_44 ;
wire un9_axb_45 ;
wire un9_6_0_cry_5_RNO ;
wire un9_6_0_cry_5 ;
wire un9_6_0_axb_6 ;
wire un9_6_0_cry_6 ;
wire un9_6_0_axb_7 ;
wire un9_6_0_cry_7 ;
wire un9_6_0_axb_8 ;
wire un9_6_0_cry_8 ;
wire un9_6_0_cry_9 ;
wire un9_6_0_axb_10 ;
wire un9_6_0_cry_10 ;
wire un9_6_0_axb_11 ;
wire un9_6_0_cry_11 ;
wire un9_6_0_axb_12 ;
wire un9_6_0_cry_12 ;
wire un9_6_0_axb_13 ;
wire un9_6_0_cry_13 ;
wire un9_6_0_axb_14 ;
wire un9_6_0_cry_14 ;
wire un9_6_0_axb_15 ;
wire un9_6_0_cry_15 ;
wire un9_6_0_axb_16 ;
wire un9_6_0_cry_16 ;
wire un9_6_0_axb_17 ;
wire un9_6_0_cry_17 ;
wire un9_6_0_axb_18 ;
wire un9_6_0_cry_18 ;
wire un9_6_0_axb_19 ;
wire un9_6_0_cry_19 ;
wire un9_6_0_axb_20 ;
wire un9_6_0_cry_20 ;
wire un9_6_0_axb_21 ;
wire un9_6_0_cry_21 ;
wire un9_6_0_axb_22 ;
wire un9_6_0_cry_22 ;
wire un9_6_0_axb_23 ;
wire un9_6_0_cry_23 ;
wire un9_6_0_axb_24 ;
wire un9_6_0_cry_24 ;
wire un9_6_0_axb_25 ;
wire un9_6_0_cry_25 ;
wire un9_6_0_axb_26 ;
wire un9_6_0_cry_26 ;
wire un9_6_0_axb_27 ;
wire un9_6_0_cry_27 ;
wire un9_6_0_axb_28 ;
wire un9_6_0_cry_28 ;
wire un9_6_0_axb_29 ;
wire un9_6_0_cry_29 ;
wire un9_6_0_cry_30_RNO ;
wire un9_6_0_axb_30 ;
wire un9_6_0_cry_30 ;
wire un9_6_0_axb_31 ;
wire un9_6_0_cry_31 ;
wire un9_6_0_cry_32_RNO ;
wire un9_6_0_axb_32 ;
wire un9_6_0_cry_32 ;
wire un9_6_0_cry_33_RNO ;
wire un9_6_0_axb_33 ;
wire un9_6_0_cry_33 ;
wire un9_6_0_cry_34_RNO ;
wire un9_6_0_axb_34 ;
wire un9_6_0_cry_34 ;
wire un9_6_0_cry_35_RNO ;
wire un9_6_0_axb_35 ;
wire un9_6_0_cry_35 ;
wire un9_6_0_cry_36_RNO ;
wire un9_6_0_axb_36 ;
wire un9_6_0_cry_36 ;
wire un9_6_0_axb_37 ;
wire un9_6_0_cry_37 ;
wire un9_6_0_axb_38 ;
wire un9_6_0_cry_38 ;
wire un9_6_0_axb_39 ;
wire un9_6_0_cry_39 ;
wire un9_6_0_axb_40 ;
wire un9_6_0_cry_40 ;
wire un9_6_0_axb_41 ;
wire un9_6_0_cry_41 ;
wire un9_6_0_axb_42 ;
wire un9_6_0_cry_42 ;
wire un9_6_0_axb_43 ;
wire un9_6_0_cry_43 ;
wire un9_6_0_axb_44 ;
wire un9_6_0_cry_44 ;
wire un9_6_0_axb_45 ;
wire un9_6_0_cry_45 ;
wire un9_6_0_axb_46 ;
wire un9_8_cry_0 ;
wire un9_8_axb_1 ;
wire un9_8_cry_1 ;
wire un9_8_axb_2 ;
wire un9_8_cry_2 ;
wire un9_8_axb_3 ;
wire un9_8_cry_3 ;
wire un9_8_axb_4 ;
wire un9_8_cry_4 ;
wire un9_8_axb_5 ;
wire un9_8_cry_5 ;
wire un9_8_cry_6_RNO ;
wire un9_8_axb_6 ;
wire un9_8_cry_6 ;
wire un9_8_axb_7 ;
wire un9_8_cry_7 ;
wire un9_8_axb_8 ;
wire un9_8_cry_8 ;
wire un9_8_axb_9 ;
wire un9_8_cry_9 ;
wire un9_8_axb_10 ;
wire un9_8_cry_10 ;
wire un9_8_axb_11 ;
wire un9_8_cry_11 ;
wire un9_8_axb_12 ;
wire un9_8_cry_12 ;
wire un9_8_axb_13 ;
wire un9_8_cry_13 ;
wire un9_8_axb_14 ;
wire un9_8_cry_14 ;
wire un9_8_axb_15 ;
wire un9_8_cry_15 ;
wire un9_8_axb_16 ;
wire un9_8_cry_16 ;
wire un9_8_axb_17 ;
wire un9_8_cry_17 ;
wire un9_8_axb_18 ;
wire un9_8_cry_18 ;
wire un9_8_axb_19 ;
wire un9_8_cry_19 ;
wire un9_8_axb_20 ;
wire un9_8_cry_20 ;
wire un9_8_axb_21 ;
wire un9_8_cry_21 ;
wire un9_8_cry_22_RNO ;
wire un9_8_axb_22 ;
wire un9_8_cry_22 ;
wire un9_8_cry_23_RNO ;
wire un9_8_axb_23 ;
wire un9_8_cry_23 ;
wire un9_8_axb_24 ;
wire un9_8_cry_24 ;
wire un9_8_axb_25 ;
wire un9_8_cry_25 ;
wire un9_8_axb_26 ;
wire un9_8_cry_26 ;
wire un9_8_axb_27 ;
wire un9_8_cry_27 ;
wire un9_8_axb_28 ;
wire un9_8_cry_28 ;
wire un9_8_axb_29 ;
wire un9_8_cry_29 ;
wire un9_8_cry_30 ;
wire un9_8_axb_31 ;
wire un9_8_cry_31 ;
wire un9_8_axb_32 ;
wire un9_8_cry_32 ;
wire un9_8_axb_33 ;
wire un9_8_cry_33 ;
wire un9_8_axb_34 ;
wire un9_8_cry_34 ;
wire un9_8_axb_35 ;
wire un9_8_axb_36 ;
wire un9_10_cry_0 ;
wire un9_10_axb_1 ;
wire un9_10_cry_1 ;
wire un9_10_axb_2 ;
wire un9_10_cry_2 ;
wire un9_10_axb_3 ;
wire un9_10_cry_3 ;
wire un9_10_cry_4_RNO ;
wire un9_10_axb_4 ;
wire un9_10_cry_4 ;
wire un9_10_cry_5_RNO ;
wire un9_10_axb_5 ;
wire un9_10_cry_5 ;
wire un9_10_axb_6 ;
wire un9_10_cry_6 ;
wire un9_10_axb_7 ;
wire un9_10_cry_7 ;
wire un9_10_cry_8_RNO ;
wire un9_10_axb_8 ;
wire un9_10_cry_8 ;
wire un9_10_axb_9 ;
wire un9_10_cry_9 ;
wire un9_10_axb_10 ;
wire un9_10_cry_10 ;
wire un9_10_axb_11 ;
wire un9_10_cry_11 ;
wire un9_10_axb_12 ;
wire un9_10_cry_12 ;
wire un9_10_axb_13 ;
wire un9_10_cry_13 ;
wire un9_10_axb_14 ;
wire un9_10_cry_14 ;
wire un9_10_axb_15 ;
wire un9_10_cry_15 ;
wire un9_10_axb_16 ;
wire un9_10_cry_16 ;
wire un9_10_axb_17 ;
wire un9_10_cry_17 ;
wire un9_10_axb_18 ;
wire un9_10_cry_18 ;
wire un9_10_axb_19 ;
wire un9_10_cry_19 ;
wire un9_10_axb_20 ;
wire un9_10_cry_20 ;
wire un9_10_axb_21 ;
wire un9_10_cry_21 ;
wire un9_10_axb_22 ;
wire un9_10_cry_22 ;
wire un9_10_axb_23 ;
wire un9_10_cry_23 ;
wire un9_10_axb_24 ;
wire un9_10_cry_24 ;
wire un9_10_cry_25_RNO ;
wire un9_10_axb_25 ;
wire un9_10_cry_25 ;
wire un9_10_cry_26_RNO ;
wire un9_10_axb_26 ;
wire un9_10_cry_26 ;
wire un9_10_cry_27_RNO ;
wire un9_10_axb_27 ;
wire un9_10_cry_27 ;
wire un9_10_axb_28 ;
wire un9_10_cry_28 ;
wire un9_10_axb_29 ;
wire un10_s_24 ;
wire un10_s_25 ;
wire un10_s_26 ;
wire un10_s_27 ;
wire un10_s_28 ;
wire un10_s_29 ;
wire un10_s_30 ;
wire un10_s_31 ;
wire un10_s_32 ;
wire un10_s_33 ;
wire un10_s_34 ;
wire un10_s_35 ;
wire un10_s_36 ;
wire un10_s_37 ;
wire un10_s_38 ;
wire un10_s_39 ;
wire un10_s_40 ;
wire un10_s_41 ;
wire un10_cry_0 ;
wire un10_axb_1 ;
wire un10_cry_1 ;
wire un10_axb_2 ;
wire un10_cry_2 ;
wire un10_axb_3 ;
wire un10_cry_3 ;
wire un10_axb_4 ;
wire un10_cry_4 ;
wire un10_axb_5 ;
wire un10_cry_5 ;
wire un10_axb_6 ;
wire un10_cry_6 ;
wire un10_axb_7 ;
wire un10_cry_7 ;
wire un10_axb_8 ;
wire un10_cry_8 ;
wire un10_axb_9 ;
wire un10_cry_9 ;
wire un10_axb_10 ;
wire un10_cry_10 ;
wire un10_axb_11 ;
wire un10_cry_11 ;
wire un10_axb_12 ;
wire un10_cry_12 ;
wire un10_axb_13 ;
wire un10_cry_13 ;
wire un10_axb_14 ;
wire un10_cry_14 ;
wire un10_axb_15 ;
wire un10_cry_15 ;
wire un10_axb_16 ;
wire un10_cry_16 ;
wire un10_axb_17 ;
wire un10_cry_17 ;
wire un10_axb_18 ;
wire un10_cry_18 ;
wire un10_axb_19 ;
wire un10_cry_19 ;
wire un10_axb_20 ;
wire un10_cry_20 ;
wire un10_axb_21 ;
wire un10_cry_21 ;
wire un10_axb_22 ;
wire un10_cry_22 ;
wire un10_axb_23 ;
wire un10_cry_23 ;
wire un10_axb_24 ;
wire un10_cry_24 ;
wire un10_axb_25 ;
wire un10_cry_25 ;
wire un10_axb_26 ;
wire un10_cry_26 ;
wire un10_axb_27 ;
wire un10_cry_27 ;
wire un10_axb_28 ;
wire un10_cry_28 ;
wire un10_axb_29 ;
wire un10_cry_29 ;
wire un10_cry_30_RNO ;
wire un10_axb_30 ;
wire un10_cry_30 ;
wire un10_axb_31 ;
wire un10_cry_31 ;
wire un10_axb_32 ;
wire un10_cry_32 ;
wire un10_axb_33 ;
wire un10_cry_33 ;
wire un10_axb_34 ;
wire un10_cry_34 ;
wire un10_axb_35 ;
wire un10_cry_35 ;
wire un10_axb_36 ;
wire un10_cry_36 ;
wire un10_axb_37 ;
wire un10_cry_37 ;
wire un10_cry_38 ;
wire un10_cry_39 ;
wire un10_cry_40 ;
wire un10_6_cry_0 ;
wire un10_6_cry_1_RNO ;
wire un10_6_axb_1 ;
wire un10_6_cry_1 ;
wire un10_6_cry_2_RNO ;
wire un10_6_axb_2 ;
wire un10_6_cry_2 ;
wire un10_6_cry_3_RNO ;
wire un10_6_axb_3 ;
wire un10_6_cry_3 ;
wire un10_6_axb_4 ;
wire un10_6_cry_4 ;
wire un10_6_axb_5 ;
wire un10_6_cry_5 ;
wire un10_6_axb_6 ;
wire un10_6_cry_6 ;
wire un10_6_axb_7 ;
wire un10_6_cry_7 ;
wire un10_6_axb_8 ;
wire un10_6_cry_8 ;
wire un10_6_axb_9 ;
wire un10_6_cry_9 ;
wire un10_6_axb_10 ;
wire un10_6_cry_10 ;
wire un10_6_axb_11 ;
wire un10_6_cry_11 ;
wire un10_6_axb_12 ;
wire un10_6_cry_12 ;
wire un10_6_axb_13 ;
wire un10_6_cry_13 ;
wire un10_6_axb_14 ;
wire un10_6_cry_14 ;
wire un10_6_axb_15 ;
wire un10_6_cry_15 ;
wire un10_6_axb_16 ;
wire un10_6_cry_16 ;
wire un10_6_axb_17 ;
wire un10_6_cry_17 ;
wire un10_6_axb_18 ;
wire un10_6_cry_18 ;
wire un10_6_axb_19 ;
wire un10_6_cry_19 ;
wire un10_6_axb_20 ;
wire un10_6_cry_20 ;
wire un10_6_cry_21_RNO ;
wire un10_6_axb_21 ;
wire un10_6_cry_21 ;
wire un10_6_cry_22_RNO ;
wire un10_6_axb_22 ;
wire un10_6_cry_22 ;
wire un10_6_cry_23_RNO ;
wire un10_6_axb_23 ;
wire un10_6_cry_23 ;
wire un10_8_34 ;
wire un10_6_axb_24 ;
wire un10_6_cry_24 ;
wire un10_8_37 ;
wire un10_6_axb_25 ;
wire un10_6_cry_25 ;
wire un10_8_40 ;
wire un10_6_axb_26 ;
wire un8_0_0_s_28 ;
wire un8_0_0_s_29 ;
wire un8_0_0_s_30 ;
wire un8_0_0_s_31 ;
wire un8_0_0_s_32 ;
wire un8_0_0_s_33 ;
wire un8_0_0_s_34 ;
wire un8_0_0_s_35 ;
wire un8_0_0_s_36 ;
wire un8_0_0_s_37 ;
wire un8_0_0_s_38 ;
wire un8_0_0_s_39 ;
wire un8_0_0_s_40 ;
wire un8_0_0_s_41 ;
wire un8_0_0_s_42 ;
wire un8_0_0_s_43 ;
wire un8_0_0_cry_0 ;
wire un8_0_0_cry_1 ;
wire un8_0_0_cry_2 ;
wire un8_0_0_cry_3 ;
wire un8_0_0_cry_4 ;
wire un8_0_0_cry_5 ;
wire un8_0_0_cry_6 ;
wire un8_0_0_axb_7 ;
wire un8_0_0_cry_7 ;
wire un8_0_0_axb_8 ;
wire un8_0_0_cry_8 ;
wire un8_0_0_axb_9 ;
wire un8_0_0_cry_9 ;
wire un8_0_0_axb_10 ;
wire un8_0_0_cry_10 ;
wire un8_0_0_axb_11 ;
wire un8_0_0_cry_11 ;
wire un8_0_0_axb_12 ;
wire un8_0_0_cry_12 ;
wire un8_0_0_axb_13 ;
wire un8_0_0_cry_13 ;
wire un8_0_0_axb_14 ;
wire un8_0_0_cry_14 ;
wire un8_0_0_axb_15 ;
wire un8_0_0_cry_15 ;
wire un8_0_0_axb_16 ;
wire un8_0_0_cry_16 ;
wire un8_0_0_axb_17 ;
wire un8_0_0_cry_17 ;
wire un8_0_0_axb_18 ;
wire un8_0_0_cry_18 ;
wire un8_0_0_axb_19 ;
wire un8_0_0_cry_19 ;
wire un8_0_0_axb_20 ;
wire un8_0_0_cry_20 ;
wire un8_0_0_axb_21 ;
wire un8_0_0_cry_21 ;
wire un8_0_0_axb_22 ;
wire un8_0_0_cry_22 ;
wire un8_0_0_axb_23 ;
wire un8_0_0_cry_23 ;
wire un8_0_0_axb_24 ;
wire un8_0_0_cry_24 ;
wire un8_0_0_axb_25 ;
wire un8_0_0_cry_25 ;
wire un8_0_0_axb_26 ;
wire un8_0_0_cry_26 ;
wire un8_0_0_axb_27 ;
wire un8_0_0_cry_27 ;
wire un8_0_0_axb_28 ;
wire un8_0_0_cry_28 ;
wire un8_0_0_axb_29 ;
wire un8_0_0_cry_29 ;
wire un8_0_0_cry_30_RNO ;
wire un8_0_0_axb_30 ;
wire un8_0_0_cry_30 ;
wire un8_0_0_cry_31_RNO ;
wire un8_0_0_axb_31 ;
wire un8_0_0_cry_31 ;
wire un8_0_0_cry_32_RNO ;
wire un8_0_0_axb_32 ;
wire un8_0_0_cry_32 ;
wire un8_0_0_cry_33_RNO ;
wire un8_0_0_axb_33 ;
wire un8_0_0_cry_33 ;
wire un8_0_0_cry_34_RNO ;
wire un8_0_0_axb_34 ;
wire un8_0_0_cry_34 ;
wire un8_0_0_cry_35_RNO ;
wire un8_0_0_axb_35 ;
wire un8_0_0_cry_35 ;
wire un8_0_0_cry_36_RNO ;
wire un8_0_0_axb_36 ;
wire un8_0_0_cry_36 ;
wire un8_0_0_axb_37 ;
wire un8_0_0_cry_37 ;
wire un8_0_0_axb_38 ;
wire un8_0_0_cry_38 ;
wire un8_0_0_axb_39 ;
wire un8_0_0_cry_39 ;
wire un8_0_0_cry_40 ;
wire un8_0_0_axb_41 ;
wire un8_0_0_cry_41 ;
wire un8_0_0_axb_42 ;
wire un8_0_0_cry_42 ;
wire un8_0_0_axb_43 ;
wire un8_0_6_cry_0 ;
wire un8_0_6_axb_1 ;
wire un8_0_6_cry_1 ;
wire un8_0_6_axb_2 ;
wire un8_0_6_cry_2 ;
wire un8_0_6_axb_3 ;
wire un8_0_6_cry_3 ;
wire un8_0_6_cry_4_RNO ;
wire un8_0_6_axb_4 ;
wire un8_0_6_cry_4 ;
wire un8_0_6_axb_5 ;
wire un8_0_6_cry_5 ;
wire un8_0_6_axb_6 ;
wire un8_0_6_cry_6 ;
wire un8_0_6_axb_7 ;
wire un8_0_6_cry_7 ;
wire un8_0_6_axb_8 ;
wire un8_0_6_cry_8 ;
wire un8_0_6_axb_9 ;
wire un8_0_6_cry_9 ;
wire un8_0_6_axb_10 ;
wire un8_0_6_cry_10 ;
wire un8_0_6_axb_11 ;
wire un8_0_6_cry_11 ;
wire un8_0_6_axb_12 ;
wire un8_0_6_cry_12 ;
wire un8_0_6_axb_13 ;
wire un8_0_6_cry_13 ;
wire un8_0_6_axb_14 ;
wire un8_0_6_cry_14 ;
wire un8_0_6_axb_15 ;
wire un8_0_6_cry_15 ;
wire un8_0_6_axb_16 ;
wire un8_0_6_cry_16 ;
wire un8_0_6_axb_17 ;
wire un8_0_6_cry_17 ;
wire un8_0_6_axb_18 ;
wire un8_0_6_cry_18 ;
wire un8_0_6_axb_19 ;
wire un8_0_6_cry_19 ;
wire un8_0_6_cry_20_RNO ;
wire un8_0_6_axb_20 ;
wire un8_0_6_cry_20 ;
wire un8_0_6_43 ;
wire un8_0_6_axb_21 ;
wire un8_0_6_cry_21 ;
wire un8_0_6_axb_22 ;
wire un7_0_0_cry_0 ;
wire un7_0_0_axb_1 ;
wire un7_0_0_cry_1 ;
wire un7_0_0_axb_2 ;
wire un7_0_0_cry_2 ;
wire un7_0_0_axb_3 ;
wire un7_0_0_cry_3 ;
wire un7_0_0_axb_4 ;
wire un7_0_0_cry_4 ;
wire un7_0_0_axb_5 ;
wire un7_0_0_cry_5 ;
wire un7_0_0_axb_6 ;
wire un7_0_0_cry_6 ;
wire un7_0_0_axb_7 ;
wire un7_0_0_cry_7 ;
wire un7_0_0_axb_8 ;
wire un7_0_0_cry_8 ;
wire un7_0_0_axb_9 ;
wire un7_0_0_cry_9 ;
wire un7_0_0_axb_10 ;
wire un7_0_0_cry_10 ;
wire un7_0_0_axb_11 ;
wire un7_0_0_cry_11 ;
wire un7_0_0_axb_12 ;
wire un7_0_0_cry_12 ;
wire un7_0_0_axb_13 ;
wire un7_0_0_cry_13 ;
wire un7_0_0_axb_14 ;
wire un7_0_0_cry_14 ;
wire un7_0_0_axb_15 ;
wire un7_0_0_cry_15 ;
wire un7_0_0_axb_16 ;
wire un7_0_0_cry_16 ;
wire un7_0_0_axb_17 ;
wire un7_0_0_cry_17 ;
wire un7_0_0_axb_18 ;
wire un7_0_0_cry_18 ;
wire un7_0_0_axb_19 ;
wire un7_0_0_cry_19 ;
wire un7_0_0_axb_20 ;
wire un7_0_0_cry_20 ;
wire un7_0_0_axb_21 ;
wire un7_0_0_cry_21 ;
wire un7_0_0_axb_22 ;
wire un7_0_0_cry_22 ;
wire un7_0_0_axb_23 ;
wire un7_0_0_cry_23 ;
wire un7_0_0_axb_24 ;
wire un7_0_0_cry_24 ;
wire un7_0_0_axb_25 ;
wire un7_0_0_cry_25 ;
wire un7_0_0_axb_26 ;
wire un7_0_0_cry_26 ;
wire un7_0_0_axb_27 ;
wire un7_0_0_cry_27 ;
wire un7_0_0_axb_28 ;
wire un7_0_0_cry_28 ;
wire un7_0_0_axb_29 ;
wire un7_0_0_cry_29 ;
wire un7_0_0_axb_30 ;
wire un7_0_0_cry_30 ;
wire un7_0_0_axb_31 ;
wire un7_0_0_cry_31 ;
wire un7_0_0_axb_32 ;
wire un7_0_0_cry_32 ;
wire un7_0_0_axb_33 ;
wire un7_0_0_cry_33 ;
wire un7_0_0_axb_34 ;
wire un7_0_0_cry_34 ;
wire un7_0_0_cry_35_RNO ;
wire un7_0_0_axb_35 ;
wire un7_0_0_cry_35 ;
wire un7_0_0_cry_36_RNO ;
wire un7_0_0_axb_36 ;
wire un7_0_0_cry_36 ;
wire un7_0_0_cry_37_RNO ;
wire un7_0_0_axb_37 ;
wire un7_0_0_cry_37 ;
wire un7_0_0_cry_38_RNO ;
wire un7_0_0_axb_38 ;
wire un7_0_0_cry_38 ;
wire un7_0_0_axb_39 ;
wire un7_0_0_cry_39 ;
wire un7_0_0_cry_40_RNO ;
wire un7_0_0_axb_40 ;
wire un7_0_0_cry_40 ;
wire un7_0_0_cry_41_RNO ;
wire un7_0_0_axb_41 ;
wire un7_0_0_cry_41 ;
wire un7_0_0_axb_42 ;
wire un7_0_0_cry_42 ;
wire un7_0_0_axb_43 ;
wire un7_0_0_cry_43 ;
wire un7_0_0_axb_44 ;
wire un7_0_0_cry_44 ;
wire un7_0_0_axb_45 ;
wire un7_0_6_cry_0 ;
wire un7_0_6_axb_1 ;
wire un7_0_6_cry_1 ;
wire un7_0_6_axb_2 ;
wire un7_0_6_cry_2 ;
wire un7_0_6_axb_3 ;
wire un7_0_6_cry_3 ;
wire un7_0_6_cry_4_RNO ;
wire un7_0_6_axb_4 ;
wire un7_0_6_cry_4 ;
wire un7_0_6_axb_5 ;
wire un7_0_6_cry_5 ;
wire un7_0_6_cry_6_RNO ;
wire un7_0_6_axb_6 ;
wire un7_0_6_cry_6 ;
wire un7_0_6_axb_7 ;
wire un7_0_6_cry_7 ;
wire un7_0_6_cry_8_RNO ;
wire un7_0_6_axb_8 ;
wire un7_0_6_cry_8 ;
wire un7_0_6_cry_9_RNO ;
wire un7_0_6_axb_9 ;
wire un7_0_6_cry_9 ;
wire un7_0_6_axb_10 ;
wire un7_0_6_cry_10 ;
wire un7_0_6_axb_11 ;
wire un7_0_6_cry_11 ;
wire un7_0_6_axb_12 ;
wire un7_0_6_cry_12 ;
wire un7_0_6_axb_13 ;
wire un7_0_6_cry_13 ;
wire un7_0_6_axb_14 ;
wire un7_0_6_cry_14 ;
wire un7_0_6_axb_15 ;
wire un7_0_6_cry_15 ;
wire un7_0_6_axb_16 ;
wire un7_0_6_cry_16 ;
wire un7_0_6_axb_17 ;
wire un7_0_6_cry_17 ;
wire un7_0_6_axb_18 ;
wire un7_0_6_cry_18 ;
wire un7_0_6_axb_19 ;
wire un7_0_6_cry_19 ;
wire un7_0_6_axb_20 ;
wire un7_0_6_cry_20 ;
wire un7_0_6_axb_21 ;
wire un7_0_6_cry_21 ;
wire un7_0_6_axb_22 ;
wire un7_0_6_cry_22 ;
wire un7_0_6_cry_23_RNO ;
wire un7_0_6_axb_23 ;
wire un7_0_6_cry_23 ;
wire un7_0_6_axb_24 ;
wire un7_0_6_cry_24 ;
wire un7_0_6_axb_25 ;
wire un7_0_6_cry_25 ;
wire un7_0_6_axb_26 ;
wire un7_0_6_cry_26 ;
wire un7_0_6_axb_27 ;
wire un7_0_6_cry_27 ;
wire un7_0_6_axb_28 ;
wire un7_0_6_cry_28 ;
wire un7_0_6_axb_29 ;
wire un7_0_8_cry_0 ;
wire un7_0_8_axb_1 ;
wire un7_0_8_cry_1 ;
wire un7_0_8_axb_2 ;
wire un7_0_8_cry_2 ;
wire un7_0_8_axb_3 ;
wire un7_0_8_cry_3 ;
wire un7_0_8_axb_4 ;
wire un7_0_8_cry_4 ;
wire un7_0_8_axb_5 ;
wire un7_0_8_cry_5 ;
wire un7_0_8_axb_6 ;
wire un7_0_8_cry_6 ;
wire un7_0_8_axb_7 ;
wire un7_0_8_cry_7 ;
wire un7_0_8_axb_8 ;
wire un7_0_8_cry_8 ;
wire un7_0_8_axb_9 ;
wire un7_0_8_cry_9 ;
wire un7_0_8_axb_10 ;
wire un7_0_8_cry_10 ;
wire un7_0_8_axb_11 ;
wire un7_0_8_cry_11 ;
wire un7_0_8_axb_12 ;
wire un7_0_8_cry_12 ;
wire un7_0_8_axb_13 ;
wire un7_0_8_cry_13 ;
wire un7_0_8_axb_14 ;
wire un7_0_8_cry_14 ;
wire un7_0_8_axb_15 ;
wire un7_0_8_cry_15 ;
wire un7_0_8_axb_16 ;
wire un7_0_8_cry_16 ;
wire un7_0_8_axb_17 ;
wire un7_0_8_cry_17 ;
wire un7_0_8_axb_18 ;
wire un7_0_8_cry_18 ;
wire un7_0_8_axb_19 ;
wire un7_0_8_cry_19 ;
wire un7_0_8_19 ;
wire un7_0_8_axb_20 ;
wire un7_0_8_cry_20 ;
wire un7_0_8_22 ;
wire un7_0_8_axb_21 ;
wire un7_0_8_cry_21 ;
wire un7_0_8_axb_22 ;
wire un7_0_8_cry_22 ;
wire un7_0_8_axb_23 ;
wire un7_0_8_cry_23 ;
wire un7_0_8_axb_24 ;
wire un7_0_8_cry_24 ;
wire un7_0_8_axb_25 ;
wire un7_0_8_cry_25 ;
wire un7_0_8_axb_26 ;
wire un7_0_8_cry_26 ;
wire un7_0_8_axb_27 ;
wire un7_0_8_cry_27 ;
wire un7_0_8_axb_28 ;
wire un6_0_8_cry_0 ;
wire un6_0_8_axb_1 ;
wire un6_0_8_cry_1 ;
wire un6_0_8_axb_2 ;
wire un6_0_8_cry_2 ;
wire un6_0_8_axb_3 ;
wire un6_0_8_cry_3 ;
wire un6_0_8_axb_4 ;
wire un6_0_8_cry_4 ;
wire un6_0_8_axb_5 ;
wire un6_0_8_cry_5 ;
wire un6_0_8_axb_6 ;
wire un6_0_8_cry_6 ;
wire un6_0_8_axb_7 ;
wire un6_0_8_cry_7 ;
wire un6_0_8_axb_8 ;
wire un6_0_8_cry_8 ;
wire un6_0_8_axb_9 ;
wire un6_0_8_cry_9 ;
wire un6_0_8_axb_10 ;
wire un6_0_8_cry_10 ;
wire un6_0_8_axb_11 ;
wire un6_0_8_cry_11 ;
wire un6_0_8_axb_12 ;
wire un6_0_8_cry_12 ;
wire un6_0_8_axb_13 ;
wire un6_0_8_cry_13 ;
wire un6_0_8_axb_14 ;
wire un6_0_8_cry_14 ;
wire un6_0_8_axb_15 ;
wire un6_0_8_cry_15 ;
wire un6_0_8_axb_16 ;
wire un6_0_8_cry_16 ;
wire un6_0_8_cry_17_RNO ;
wire un6_0_8_axb_17 ;
wire un6_0_8_cry_17 ;
wire un6_0_8_axb_18 ;
wire un6_0_8_cry_18 ;
wire un6_0_8_cry_19_RNO ;
wire un6_0_8_axb_19 ;
wire un6_0_8_cry_19 ;
wire un6_0_8_axb_20 ;
wire un6_0_8_cry_20 ;
wire un6_0_8_axb_21 ;
wire un6_0_8_cry_21 ;
wire un6_0_8_axb_22 ;
wire un6_0_8_cry_22 ;
wire un6_0_8_axb_23 ;
wire un6_0_8_cry_23 ;
wire un6_0_8_axb_24 ;
wire un6_0_8_cry_24 ;
wire un6_0_8_axb_25 ;
wire un6_0_8_cry_25 ;
wire un6_0_8_axb_26 ;
wire un6_0_8_axb_27 ;
wire un8_0_8_cry_0 ;
wire un8_0_8_axb_1 ;
wire un8_0_8_cry_1 ;
wire un8_0_8_axb_2 ;
wire un8_0_8_cry_2 ;
wire un8_0_8_axb_3 ;
wire un8_0_8_cry_3 ;
wire un8_0_8_axb_4 ;
wire un8_0_8_cry_4 ;
wire un8_0_8_axb_5 ;
wire un8_0_8_cry_5 ;
wire un8_0_8_axb_6 ;
wire un8_0_8_cry_6 ;
wire un8_0_8_axb_7 ;
wire un8_0_8_cry_7 ;
wire un8_0_8_axb_8 ;
wire un8_0_8_cry_8 ;
wire un8_0_8_axb_9 ;
wire un8_0_8_cry_9 ;
wire un8_0_8_axb_10 ;
wire un8_0_8_cry_10 ;
wire un8_0_8_axb_11 ;
wire un8_0_8_cry_11 ;
wire un8_0_8_axb_12 ;
wire un8_0_8_cry_12 ;
wire un8_0_8_axb_13 ;
wire un8_0_8_cry_13 ;
wire un8_0_8_axb_14 ;
wire un8_0_8_cry_14 ;
wire un8_0_8_axb_15 ;
wire un8_0_8_cry_15 ;
wire un8_0_8_axb_16 ;
wire un8_0_8_cry_16 ;
wire un8_0_8_cry_17_RNO ;
wire un8_0_8_axb_17 ;
wire un8_0_8_cry_17 ;
wire un8_0_8_axb_18 ;
wire un8_0_8_cry_18 ;
wire un8_0_8_cry_19_RNO ;
wire un8_0_8_axb_19 ;
wire un8_0_8_cry_19 ;
wire un8_0_8_axb_20 ;
wire un8_0_8_cry_20 ;
wire un8_0_8_axb_21 ;
wire un8_0_8_cry_21 ;
wire un8_0_8_axb_22 ;
wire un8_0_8_cry_22 ;
wire un8_0_8_axb_23 ;
wire un8_0_8_cry_23 ;
wire un8_0_8_axb_24 ;
wire un8_0_8_cry_24 ;
wire un8_0_8_axb_25 ;
wire un8_0_8_cry_25 ;
wire un8_0_8_axb_26 ;
wire un8_0_8_axb_27 ;
wire un10_8_axb_0 ;
wire un10_8_cry_0 ;
wire un10_8_axb_1 ;
wire un10_8_cry_1 ;
wire un10_8_axb_2 ;
wire un10_8_cry_2 ;
wire un10_8_axb_3 ;
wire un10_8_cry_3 ;
wire un10_8_axb_4 ;
wire un10_8_cry_4 ;
wire un10_8_axb_5 ;
wire un10_8_cry_5 ;
wire un10_8_axb_6 ;
wire un10_8_cry_6 ;
wire un10_8_axb_7 ;
wire un10_8_cry_7 ;
wire un10_8_axb_8 ;
wire un10_8_cry_8 ;
wire un10_8_axb_9 ;
wire un10_8_cry_9 ;
wire un10_8_axb_10 ;
wire un10_8_cry_10 ;
wire un10_8_cry_11_RNO ;
wire un10_8_axb_11 ;
wire un10_8_cry_11 ;
wire un10_8_axb_12 ;
wire un10_8_cry_12 ;
wire un10_8_axb_13 ;
wire un10_8_cry_13 ;
wire un10_8_axb_14 ;
wire un10_8_cry_14 ;
wire un10_8_axb_15 ;
wire un10_8_cry_15 ;
wire un10_8_axb_16 ;
wire un10_8_cry_16 ;
wire un10_8_axb_17 ;
wire un10_8_cry_17 ;
wire un10_8_axb_18 ;
wire un10_8_cry_18 ;
wire un10_8_axb_19 ;
wire un10_8_cry_19 ;
wire un10_8_axb_20 ;
wire un10_8_cry_20 ;
wire un10_8_axb_21 ;
wire un10_8_cry_21 ;
wire un10_8_axb_22 ;
wire un10_8_cry_22 ;
wire un10_8_axb_23 ;
wire un10_8_cry_23 ;
wire un10_8_axb_24 ;
wire un10_8_cry_24 ;
wire un10_8_axb_25 ;
wire un10_8_cry_25 ;
wire un10_8_axb_26 ;
wire un10_8_cry_26 ;
wire un10_8_axb_27 ;
wire un10_8_cry_27 ;
wire un10_8_axb_28 ;
wire Y_out_double_2_cry_0 ;
wire Y_out_double_2_axb_1 ;
wire Y_out_double_2_cry_1 ;
wire Y_out_double_2_axb_2 ;
wire Y_out_double_2_cry_2 ;
wire Y_out_double_2_axb_3 ;
wire Y_out_double_2_cry_3 ;
wire Y_out_double_2_axb_4 ;
wire Y_out_double_2_cry_4 ;
wire Y_out_double_2_axb_5 ;
wire Y_out_double_2_cry_5 ;
wire Y_out_double_2_axb_6 ;
wire Y_out_double_2_cry_6 ;
wire Y_out_double_2_axb_7 ;
wire Y_out_double_2_cry_7 ;
wire Y_out_double_2_axb_8 ;
wire Y_out_double_2_cry_8 ;
wire Y_out_double_2_axb_9 ;
wire Y_out_double_2_cry_9 ;
wire Y_out_double_2_axb_10 ;
wire Y_out_double_2_cry_10 ;
wire Y_out_double_2_axb_11 ;
wire Y_out_double_2_cry_11 ;
wire Y_out_double_2_axb_12 ;
wire Y_out_double_2_cry_12 ;
wire Y_out_double_2_axb_13 ;
wire Y_out_double_2_cry_13 ;
wire Y_out_double_2_axb_14 ;
wire Y_out_double_2_cry_14 ;
wire Y_out_double_2_axb_15 ;
wire Y_out_double_2_cry_15 ;
wire Y_out_double_2_axb_16 ;
wire Y_out_double_2_cry_16 ;
wire Y_out_double_2_axb_17 ;
wire Y_out_double_2_7_cry_1 ;
wire Y_out_double_2_7_axb_2 ;
wire Y_out_double_2_7_cry_2 ;
wire Y_out_double_2_7_axb_3 ;
wire Y_out_double_2_7_cry_3 ;
wire Y_out_double_2_7_axb_4 ;
wire Y_out_double_2_7_cry_4 ;
wire Y_out_double_2_7_axb_5 ;
wire Y_out_double_2_7_cry_5 ;
wire Y_out_double_2_7_axb_6 ;
wire Y_out_double_2_7_cry_6 ;
wire Y_out_double_2_7_axb_7 ;
wire Y_out_double_2_7_cry_7 ;
wire Y_out_double_2_7_axb_8 ;
wire Y_out_double_2_7_cry_8 ;
wire Y_out_double_2_7_axb_9 ;
wire Y_out_double_2_7_cry_9 ;
wire Y_out_double_2_7_axb_10 ;
wire Y_out_double_2_7_cry_10 ;
wire Y_out_double_2_7_axb_11 ;
wire Y_out_double_2_7_cry_11 ;
wire Y_out_double_2_7_axb_12 ;
wire Y_out_double_2_7_cry_12 ;
wire Y_out_double_2_7_axb_13 ;
wire Y_out_double_2_7_cry_13 ;
wire Y_out_double_2_7_axb_14 ;
wire Y_out_double_2_7_cry_14 ;
wire Y_out_double_2_7_axb_15 ;
wire Y_out_double_2_7_cry_15 ;
wire Y_out_double_2_7_axb_16 ;
wire un6_0_9_cry_0 ;
wire un6_0_9_axb_1 ;
wire un6_0_9_cry_1 ;
wire un6_0_9_axb_2 ;
wire un6_0_9_cry_2 ;
wire un6_0_9_axb_3 ;
wire un6_0_9_cry_3 ;
wire un6_0_9_axb_4 ;
wire un6_0_9_cry_4 ;
wire un6_0_9_axb_5 ;
wire un6_0_9_cry_5 ;
wire un6_0_9_axb_6 ;
wire un6_0_9_cry_6 ;
wire un6_0_9_axb_7 ;
wire un6_0_9_cry_7 ;
wire un6_0_9_axb_8 ;
wire un6_0_9_cry_8 ;
wire un6_0_9_axb_9 ;
wire un6_0_9_cry_9 ;
wire un6_0_9_axb_10 ;
wire un6_0_9_cry_10 ;
wire un6_0_9_axb_11 ;
wire un6_0_9_cry_11 ;
wire un6_0_9_axb_12 ;
wire un6_0_9_cry_12 ;
wire un6_0_9_axb_13 ;
wire un6_0_9_cry_13 ;
wire un6_0_9_axb_14 ;
wire un6_0_9_cry_14 ;
wire un6_0_9_axb_15 ;
wire un6_0_9_cry_15 ;
wire un6_0_9_axb_16 ;
wire un6_0_9_cry_16 ;
wire un6_0_9_axb_17 ;
wire un6_0_9_cry_17 ;
wire un6_0_9_axb_18 ;
wire un6_0_9_cry_18 ;
wire un6_0_9_axb_19 ;
wire un6_0_9_cry_19 ;
wire un6_0_9_axb_20 ;
wire un6_0_9_cry_20 ;
wire un6_0_9_axb_21 ;
wire un6_0_9_cry_21 ;
wire un6_0_9_axb_22 ;
wire un6_0_9_cry_22 ;
wire un6_0_9_axb_23 ;
wire un6_0_9_cry_23 ;
wire un6_0_9_axb_24 ;
wire un6_0_9_cry_24 ;
wire un6_0_9_axb_25 ;
wire un6_0_9_cry_25 ;
wire un6_0_9_axb_26 ;
wire un8_0_9_cry_0 ;
wire un8_0_9_axb_1 ;
wire un8_0_9_cry_1 ;
wire un8_0_9_axb_2 ;
wire un8_0_9_cry_2 ;
wire un8_0_9_axb_3 ;
wire un8_0_9_cry_3 ;
wire un8_0_9_axb_4 ;
wire un8_0_9_cry_4 ;
wire un8_0_9_axb_5 ;
wire un8_0_9_cry_5 ;
wire un8_0_9_axb_6 ;
wire un8_0_9_cry_6 ;
wire un8_0_9_axb_7 ;
wire un8_0_9_cry_7 ;
wire un8_0_9_axb_8 ;
wire un8_0_9_cry_8 ;
wire un8_0_9_axb_9 ;
wire un8_0_9_cry_9 ;
wire un8_0_9_axb_10 ;
wire un8_0_9_cry_10 ;
wire un8_0_9_axb_11 ;
wire un8_0_9_cry_11 ;
wire un8_0_9_axb_12 ;
wire un8_0_9_cry_12 ;
wire un8_0_9_axb_13 ;
wire un8_0_9_cry_13 ;
wire un8_0_9_axb_14 ;
wire un8_0_9_cry_14 ;
wire un8_0_9_axb_15 ;
wire un8_0_9_cry_15 ;
wire un8_0_9_axb_16 ;
wire un8_0_9_cry_16 ;
wire un8_0_9_axb_17 ;
wire un8_0_9_cry_17 ;
wire un8_0_9_axb_18 ;
wire un8_0_9_cry_18 ;
wire un8_0_9_axb_19 ;
wire un8_0_9_cry_19 ;
wire un8_0_9_axb_20 ;
wire un8_0_9_cry_20 ;
wire un8_0_9_axb_21 ;
wire un8_0_9_cry_21 ;
wire un8_0_9_axb_22 ;
wire un8_0_9_cry_22 ;
wire un8_0_9_axb_23 ;
wire un8_0_9_cry_23 ;
wire un8_0_9_axb_24 ;
wire un8_0_9_cry_24 ;
wire un8_0_9_axb_25 ;
wire un8_0_9_cry_25 ;
wire un8_0_9_axb_26 ;
wire un9_11_cry_6 ;
wire un9_11_axb_7 ;
wire un9_11_cry_7 ;
wire un9_11_axb_8 ;
wire un9_11_cry_8 ;
wire un9_11_axb_9 ;
wire un9_11_cry_9 ;
wire un9_11_axb_10 ;
wire un9_11_cry_10 ;
wire un9_11_axb_11 ;
wire un9_11_cry_11 ;
wire un9_11_axb_12 ;
wire un9_11_cry_12 ;
wire un9_11_axb_13 ;
wire un9_11_cry_13 ;
wire un9_11_axb_14 ;
wire un9_11_cry_14 ;
wire un9_11_axb_15 ;
wire un9_11_cry_15 ;
wire un9_11_axb_16 ;
wire un9_11_cry_16 ;
wire un9_11_axb_17 ;
wire un9_11_cry_17 ;
wire un9_11_axb_18 ;
wire un9_11_cry_18 ;
wire un9_11_axb_19 ;
wire un9_11_cry_19 ;
wire un9_11_axb_20 ;
wire un9_11_cry_20 ;
wire un9_11_axb_21 ;
wire un9_11_cry_21 ;
wire un9_11_axb_22 ;
wire un9_11_cry_22 ;
wire un9_11_axb_23 ;
wire un9_11_cry_23 ;
wire un9_11_axb_24 ;
wire Y_out_double_2_4_cry_0 ;
wire Y_out_double_2_4_axb_1 ;
wire Y_out_double_2_4_cry_1 ;
wire Y_out_double_2_4_axb_2 ;
wire Y_out_double_2_4_cry_2 ;
wire Y_out_double_2_4_axb_3 ;
wire Y_out_double_2_4_cry_3 ;
wire Y_out_double_2_4_axb_4 ;
wire Y_out_double_2_4_cry_4 ;
wire Y_out_double_2_4_axb_5 ;
wire Y_out_double_2_4_cry_5 ;
wire Y_out_double_2_4_axb_6 ;
wire Y_out_double_2_4_cry_6 ;
wire Y_out_double_2_4_axb_7 ;
wire Y_out_double_2_4_cry_7 ;
wire Y_out_double_2_4_axb_8 ;
wire Y_out_double_2_4_cry_8 ;
wire Y_out_double_2_4_axb_9 ;
wire Y_out_double_2_4_cry_9 ;
wire Y_out_double_2_4_axb_10 ;
wire Y_out_double_2_4_cry_10 ;
wire Y_out_double_2_4_axb_11 ;
wire Y_out_double_2_4_cry_11 ;
wire Y_out_double_2_4_axb_12 ;
wire Y_out_double_2_4_cry_12 ;
wire Y_out_double_2_4_axb_13 ;
wire Y_out_double_2_4_cry_13 ;
wire Y_out_double_2_4_axb_14 ;
wire Y_out_double_2_4_cry_14 ;
wire Y_out_double_2_4_axb_15 ;
wire Y_out_double_2_4_cry_15 ;
wire Y_out_double_2_4_axb_16 ;
wire Y_out_double_2_4_cry_16 ;
wire Y_out_double_2_4_axb_17 ;
wire N_2197_i ;
wire N_2393_i ;
wire N_3207_i ;
wire N_3204_i ;
wire N_3201_i ;
wire N_3198_i ;
wire N_3195_i ;
wire N_3193_i ;
wire N_3186_i ;
wire N_2390_i ;
wire N_2387_i ;
wire N_2384_i ;
wire N_2381_i ;
wire N_2379_i ;
wire N_2372_i ;
wire N_3387_i ;
wire N_3385_i ;
wire N_3180_i ;
wire N_1128_i ;
wire N_2973_i ;
wire N_2366_i ;
wire N_2007_i ;
wire N_3313_i ;
wire n_reset_i ;
wire un8_0_0_cry_6_sf ;
wire un10_cry_40_sf ;
wire un6_0_0_cry_6_sf ;
wire un8_0_6_cry_0_sf ;
wire un6_0_6_cry_0_sf ;
wire un9_11_cry_6_RNO ;
wire un10_6_cry_0_RNO_0 ;
wire un9_8_cry_30_RNO ;
wire un9_8_cry_0_RNO ;
wire un9_6_0_cry_9_RNO ;
wire un9_6_0_cry_5_RNO_0 ;
wire un10_8_cry_0_cy ;
wire un9_cry_0_cy ;
wire un9_10_8_rep1 ;
wire ZFF_Y1_15_rep1 ;
wire ZFF_X0_7_rep1 ;
wire ZFF_Y1_16_rep1 ;
wire ZFF_X0_6_rep1 ;
wire un9_8_7_rep1 ;
wire ZFF_X0_10_rep1 ;
wire ZFF_X0_11_rep1 ;
wire ZFF_X0_12_rep1 ;
wire ZFF_X2_6_rep1 ;
wire ZFF_X0_4_rep1 ;
wire ZFF_X2_10_rep1 ;
wire ZFF_X0_2_rep1 ;
wire ZFF_X0_1_rep1 ;
wire un9_8_6_rep1 ;
wire ZFF_X2_2_rep1 ;
wire ZFF_X0_3_rep1 ;
wire ZFF_X2_3_rep1 ;
wire ZFF_Y1_4_rep1 ;
wire ZFF_Y1_3_rep1 ;
wire ZFF_Y1_5_rep1 ;
wire ZFF_X2_14_rep1 ;
wire ZFF_X0_14_rep1 ;
wire ZFF_X0_15_rep1 ;
wire ZFF_X2_15_rep1 ;
wire ZFF_Y1_6_rep1 ;
wire un9_11_25_rep1 ;
wire ZFF_Y1_7_rep1 ;
wire un9_11_26_rep1 ;
wire ZFF_X1_3_rep1 ;
wire ZFF_X1_0_rep1 ;
wire ZFF_Y1_9_rep1 ;
wire ZFF_X1_7_rep1 ;
wire ZFF_X1_4_rep1 ;
wire ZFF_X1_1_rep1 ;
wire un9_11_22_rep1 ;
wire ZFF_X1_8_rep1 ;
wire ZFF_X1_9_rep1 ;
wire ZFF_X1_11_rep1 ;
wire ZFF_X1_15_rep1 ;
wire ZFF_X1_2_rep1 ;
wire un9_11_24_rep1 ;
wire ZFF_X0_16_rep1 ;
wire ZFF_Y1_17_rep1 ;
wire ZFF_X1_5_rep1 ;
wire ZFF_Y1_8_rep1 ;
wire ZFF_X1_6_rep1 ;
wire ZFF_X1_12_rep1 ;
wire ZFF_X1_10_rep1 ;
wire ZFF_X1_13_rep1 ;
wire un9_11_23_rep1 ;
wire ZFF_Y2_8_rep1 ;
wire ZFF_Y2_6_rep1 ;
wire ZFF_Y2_7_rep1 ;
wire ZFF_Y2_14_rep1 ;
wire un8_0_0_axb_42_N_2L1 ;
wire un6_0_0_axb_42_N_2L1 ;
wire N_3353_i_0 ;
wire un9_8_cry_29_0 ;
wire un9_8_cry_29_1 ;
wire un9_6_0_cry_8_0 ;
wire un9_6_0_cry_8_1 ;
wire un7_0_10_s_27_true ;
input p_desc86_p_O_FDE ;
input p_desc87_p_O_FDE ;
input p_desc88_p_O_FDE ;
input p_desc89_p_O_FDE ;
input p_desc90_p_O_FDE ;
input p_desc91_p_O_FDE ;
input p_desc92_p_O_FDE ;
input p_desc93_p_O_FDE ;
input p_desc94_p_O_FDE ;
input p_desc95_p_O_FDE ;
input p_desc96_p_O_FDE ;
input p_desc97_p_O_FDE ;
input p_desc98_p_O_FDE ;
input p_desc99_p_O_FDE ;
input p_desc100_p_O_FDE ;
input p_desc101_p_O_FDE ;
input p_desc102_p_O_FDE ;
input p_desc103_p_O_FDE ;
input p_desc104_p_O_FDE ;
input p_desc105_p_O_FDE ;
input p_desc106_p_O_FDE ;
input p_desc107_p_O_FDE ;
input p_desc108_p_O_FDE ;
input p_desc109_p_O_FDE ;
input p_desc110_p_O_FDE ;
input p_desc111_p_O_FDE ;
input p_desc112_p_O_FDE ;
input p_desc113_p_O_FDE ;
input p_desc114_p_O_FDE ;
input p_desc115_p_O_FDE ;
input p_desc116_p_O_FDE ;
input p_desc117_p_O_FDE ;
input p_desc118_p_O_FDE ;
input p_desc119_p_O_FDE ;
input p_desc120_p_O_FDE ;
input p_desc121_p_O_FDE ;
input p_desc162_p_O_FDE ;
input p_desc163_p_O_FDE ;
input p_desc164_p_O_FDE ;
input p_desc165_p_O_FDE ;
input p_desc166_p_O_FDE ;
input p_desc167_p_O_FDE ;
input p_desc168_p_O_FDE ;
input p_desc169_p_O_FDE ;
input p_desc170_p_O_FDE ;
input p_desc171_p_O_FDE ;
input p_desc172_p_O_FDE ;
input p_desc173_p_O_FDE ;
input p_desc174_p_O_FDE ;
input p_desc175_p_O_FDE ;
input p_desc176_p_O_FDE ;
input p_desc177_p_O_FDE ;
input p_desc178_p_O_FDE ;
input p_desc179_p_O_FDE ;
input p_desc198_p_O_FDE ;
input p_desc199_p_O_FDE ;
input p_desc200_p_O_FDE ;
input p_desc201_p_O_FDE ;
input p_desc202_p_O_FDE ;
input p_desc203_p_O_FDE ;
input p_desc204_p_O_FDE ;
input p_desc205_p_O_FDE ;
input p_desc206_p_O_FDE ;
input p_desc207_p_O_FDE ;
input p_desc208_p_O_FDE ;
input p_desc209_p_O_FDE ;
input p_desc210_p_O_FDE ;
input p_desc211_p_O_FDE ;
input p_desc212_p_O_FDE ;
input p_desc213_p_O_FDE ;
input p_desc214_p_O_FDE ;
input p_desc215_p_O_FDE ;
input p_desc216_p_O_FDE ;
input p_desc217_p_O_FDE ;
input p_desc218_p_O_FDE ;
input p_desc219_p_O_FDE ;
input p_desc220_p_O_FDE ;
input p_desc221_p_O_FDE ;
input p_desc222_p_O_FDE ;
input p_desc223_p_O_FDE ;
input p_desc224_p_O_FDE ;
input p_desc225_p_O_FDE ;
input p_desc226_p_O_FDE ;
input p_desc227_p_O_FDE ;
input p_desc228_p_O_FDE ;
input p_desc229_p_O_FDE ;
input p_desc230_p_O_FDE ;
input p_desc231_p_O_FDE ;
input p_desc232_p_O_FDE ;
input p_desc233_p_O_FDE ;
input p_desc234_p_O_FDE ;
input p_desc235_p_O_FDE ;
input p_desc236_p_O_FDE ;
input p_desc237_p_O_FDE ;
input p_desc238_p_O_FDE ;
input p_desc239_p_O_FDE ;
input p_desc240_p_O_FDE ;
input p_desc241_p_O_FDE ;
input p_desc242_p_O_FDE ;
input p_desc243_p_O_FDE ;
input p_desc244_p_O_FDE ;
input p_desc245_p_O_FDE ;
input p_desc246_p_O_FDE ;
input p_desc247_p_O_FDE ;
input p_desc248_p_O_FDE ;
input p_desc249_p_O_FDE ;
input p_desc250_p_O_FDE ;
input p_desc251_p_O_FDE ;
input p_desc252_p_O_FDE ;
input p_desc253_p_O_FDE ;
input p_desc254_p_O_FDE ;
input p_desc255_p_O_FDE ;
input p_desc256_p_O_FDE ;
input p_desc257_p_O_FDE ;
input p_desc258_p_O_FDE ;
input p_desc259_p_O_FDE ;
input p_desc260_p_O_FDE ;
input p_desc261_p_O_FDE ;
input p_desc262_p_O_FDE ;
input p_desc263_p_O_FDE ;
input p_desc264_p_O_FDE ;
input p_desc334_p_O_FDC ;
input p_desc335_p_O_FDC ;
input p_desc336_p_O_FDC ;
input p_desc337_p_O_FDC ;
input p_state_reg_ret_5_Z_p_O_FDC ;
input p_state_reg_ret_Z_p_O_FDP ;
input p_state_reg_ret_1_Z_p_O_FDP ;
input p_state_reg_ret_2_Z_p_O_FDP ;
input p_state_reg_ret_4_Z_p_O_FDP ;
input p_desc180_p_O_FDCE ;
input p_desc181_p_O_FDCE ;
input p_desc182_p_O_FDCE ;
input p_desc183_p_O_FDCE ;
input p_desc184_p_O_FDCE ;
input p_desc185_p_O_FDCE ;
input p_desc186_p_O_FDCE ;
input p_desc187_p_O_FDCE ;
input p_desc188_p_O_FDCE ;
input p_desc189_p_O_FDCE ;
input p_desc190_p_O_FDCE ;
input p_desc191_p_O_FDCE ;
input p_desc192_p_O_FDCE ;
input p_desc193_p_O_FDCE ;
input p_desc194_p_O_FDCE ;
input p_desc195_p_O_FDCE ;
input p_desc196_p_O_FDCE ;
input p_desc197_p_O_FDCE ;
input p_desc265_p_O_FDCE ;
input p_desc266_p_O_FDCE ;
input p_desc267_p_O_FDCE ;
input p_desc268_p_O_FDCE ;
input p_desc269_p_O_FDCE ;
input p_desc270_p_O_FDCE ;
input p_desc271_p_O_FDCE ;
input p_desc272_p_O_FDCE ;
input p_desc273_p_O_FDCE ;
input p_desc274_p_O_FDCE ;
input p_desc275_p_O_FDCE ;
input p_desc276_p_O_FDCE ;
input p_desc277_p_O_FDCE ;
input p_desc278_p_O_FDCE ;
input p_desc279_p_O_FDCE ;
input p_desc280_p_O_FDCE ;
input p_desc281_p_O_FDCE ;
input p_desc282_p_O_FDCE ;
input p_desc283_p_O_FDCE ;
input p_desc284_p_O_FDCE ;
input p_desc285_p_O_FDCE ;
input p_desc286_p_O_FDCE ;
input p_desc287_p_O_FDCE ;
input p_desc288_p_O_FDCE ;
input p_desc289_p_O_FDCE ;
input p_desc290_p_O_FDCE ;
input p_desc291_p_O_FDCE ;
input p_desc292_p_O_FDCE ;
input p_desc293_p_O_FDCE ;
input p_desc294_p_O_FDCE ;
input p_desc295_p_O_FDCE ;
input p_desc296_p_O_FDCE ;
input p_desc297_p_O_FDCE ;
input p_desc298_p_O_FDCE ;
input p_desc299_p_O_FDCE ;
input p_desc300_p_O_FDCE ;
input p_desc301_p_O_FDCE ;
input p_desc302_p_O_FDCE ;
input p_desc303_p_O_FDCE ;
input p_desc304_p_O_FDCE ;
input p_desc305_p_O_FDCE ;
input p_desc306_p_O_FDCE ;
input p_desc307_p_O_FDCE ;
input p_desc308_p_O_FDCE ;
input p_desc309_p_O_FDCE ;
input p_desc310_p_O_FDCE ;
input p_desc311_p_O_FDCE ;
input p_desc312_p_O_FDCE ;
input p_desc313_p_O_FDCE ;
input p_desc314_p_O_FDCE ;
input p_desc315_p_O_FDCE ;
input p_desc316_p_O_FDCE ;
input p_desc317_p_O_FDCE ;
input p_desc318_p_O_FDCE ;
input p_desc319_p_O_FDCE ;
input p_desc320_p_O_FDCE ;
input p_desc321_p_O_FDCE ;
input p_desc322_p_O_FDCE ;
input p_desc323_p_O_FDCE ;
input p_desc324_p_O_FDCE ;
input p_desc325_p_O_FDCE ;
input p_desc326_p_O_FDCE ;
input p_desc327_p_O_FDCE ;
input p_desc328_p_O_FDCE ;
input p_desc329_p_O_FDCE ;
input p_desc330_p_O_FDCE ;
input p_desc331_p_O_FDCE ;
input p_desc332_p_O_FDCE ;
input p_desc333_p_O_FDCE ;
input p_desc338_p_O_FDCE ;
input p_ZFF_Y1_0_rep1_Z_p_O_FDCE ;
input p_desc339_p_O_FDCE ;
input p_ZFF_Y1_15_rep1_Z_p_O_FDCE ;
input p_desc340_p_O_FDCE ;
input p_ZFF_X0_7_rep1_Z_p_O_FDCE ;
input p_desc341_p_O_FDCE ;
input p_desc342_p_O_FDCE ;
input p_desc343_p_O_FDCE ;
input p_desc344_p_O_FDCE ;
input p_ZFF_Y1_16_rep1_Z_p_O_FDCE ;
input p_desc345_p_O_FDCE ;
input p_ZFF_X0_6_rep1_Z_p_O_FDCE ;
input p_desc346_p_O_FDCE ;
input p_desc347_p_O_FDCE ;
input p_ZFF_Y1_2_rep1_Z_p_O_FDCE ;
input p_desc348_p_O_FDCE ;
input p_desc349_p_O_FDCE ;
input p_ZFF_X0_10_rep1_Z_p_O_FDCE ;
input p_desc350_p_O_FDCE ;
input p_ZFF_X0_11_rep1_Z_p_O_FDCE ;
input p_desc351_p_O_FDCE ;
input p_ZFF_X0_12_rep1_Z_p_O_FDCE ;
input p_desc352_p_O_FDCE ;
input p_ZFF_X2_6_rep1_Z_p_O_FDCE ;
input p_desc353_p_O_FDCE ;
input p_ZFF_X0_4_rep1_Z_p_O_FDCE ;
input p_desc354_p_O_FDCE ;
input p_desc355_p_O_FDCE ;
input p_desc356_p_O_FDCE ;
input p_desc357_p_O_FDCE ;
input p_ZFF_X2_10_rep1_Z_p_O_FDCE ;
input p_desc358_p_O_FDCE ;
input p_ZFF_X0_2_rep1_Z_p_O_FDCE ;
input p_desc359_p_O_FDCE ;
input p_ZFF_X0_1_rep1_Z_p_O_FDCE ;
input p_desc360_p_O_FDCE ;
input p_ZFF_Y1_1_rep1_Z_p_O_FDCE ;
input p_desc361_p_O_FDCE ;
input p_desc362_p_O_FDCE ;
input p_desc363_p_O_FDCE ;
input p_desc364_p_O_FDCE ;
input p_ZFF_X2_2_rep1_Z_p_O_FDCE ;
input p_desc365_p_O_FDCE ;
input p_ZFF_X0_3_rep1_Z_p_O_FDCE ;
input p_desc366_p_O_FDCE ;
input p_desc367_p_O_FDCE ;
input p_ZFF_X2_3_rep1_Z_p_O_FDCE ;
input p_desc368_p_O_FDCE ;
input p_ZFF_Y1_4_rep1_Z_p_O_FDCE ;
input p_desc369_p_O_FDCE ;
input p_desc370_p_O_FDCE ;
input p_ZFF_Y1_3_rep1_Z_p_O_FDCE ;
input p_desc371_p_O_FDCE ;
input p_desc372_p_O_FDCE ;
input p_desc373_p_O_FDCE ;
input p_ZFF_Y1_5_rep1_Z_p_O_FDCE ;
input p_desc374_p_O_FDCE ;
input p_ZFF_X2_14_rep1_Z_p_O_FDCE ;
input p_desc375_p_O_FDCE ;
input p_ZFF_X0_14_rep1_Z_p_O_FDCE ;
input p_desc376_p_O_FDCE ;
input p_ZFF_X0_15_rep1_Z_p_O_FDCE ;
input p_desc377_p_O_FDCE ;
input p_ZFF_X2_15_rep1_Z_p_O_FDCE ;
input p_desc378_p_O_FDCE ;
input p_ZFF_Y1_6_rep1_Z_p_O_FDCE ;
input p_desc379_p_O_FDCE ;
input p_ZFF_Y1_13_rep1_Z_p_O_FDCE ;
input p_desc380_p_O_FDCE ;
input p_ZFF_Y1_7_rep1_Z_p_O_FDCE ;
input p_desc381_p_O_FDCE ;
input p_ZFF_Y1_14_rep1_Z_p_O_FDCE ;
input p_desc382_p_O_FDCE ;
input p_ZFF_X1_3_rep1_Z_p_O_FDCE ;
input p_desc383_p_O_FDCE ;
input p_ZFF_X1_0_rep1_Z_p_O_FDCE ;
input p_desc384_p_O_FDCE ;
input p_ZFF_Y1_9_rep1_Z_p_O_FDCE ;
input p_desc385_p_O_FDCE ;
input p_ZFF_X1_7_rep1_Z_p_O_FDCE ;
input p_desc386_p_O_FDCE ;
input p_ZFF_X1_4_rep1_Z_p_O_FDCE ;
input p_desc387_p_O_FDCE ;
input p_ZFF_X1_1_rep1_Z_p_O_FDCE ;
input p_desc388_p_O_FDCE ;
input p_ZFF_Y1_10_rep1_Z_p_O_FDCE ;
input p_desc389_p_O_FDCE ;
input p_ZFF_X1_8_rep1_Z_p_O_FDCE ;
input p_desc390_p_O_FDCE ;
input p_ZFF_X1_9_rep1_Z_p_O_FDCE ;
input p_desc391_p_O_FDCE ;
input p_ZFF_X1_11_rep1_Z_p_O_FDCE ;
input p_desc392_p_O_FDCE ;
input p_ZFF_X1_15_rep1_Z_p_O_FDCE ;
input p_desc393_p_O_FDCE ;
input p_ZFF_X1_2_rep1_Z_p_O_FDCE ;
input p_desc394_p_O_FDCE ;
input p_ZFF_Y1_12_rep1_Z_p_O_FDCE ;
input p_desc395_p_O_FDCE ;
input p_ZFF_X0_16_rep1_Z_p_O_FDCE ;
input p_desc396_p_O_FDCE ;
input p_desc397_p_O_FDCE ;
input p_ZFF_Y1_17_rep1_Z_p_O_FDCE ;
input p_desc398_p_O_FDCE ;
input p_ZFF_X1_5_rep1_Z_p_O_FDCE ;
input p_desc399_p_O_FDCE ;
input p_ZFF_Y1_8_rep1_Z_p_O_FDCE ;
input p_desc400_p_O_FDCE ;
input p_desc401_p_O_FDCE ;
input p_desc402_p_O_FDCE ;
input p_ZFF_X1_6_rep1_Z_p_O_FDCE ;
input p_desc403_p_O_FDCE ;
input p_ZFF_X1_12_rep1_Z_p_O_FDCE ;
input p_desc404_p_O_FDCE ;
input p_ZFF_X1_10_rep1_Z_p_O_FDCE ;
input p_desc405_p_O_FDCE ;
input p_ZFF_X1_13_rep1_Z_p_O_FDCE ;
input p_desc406_p_O_FDCE ;
input p_ZFF_Y1_11_rep1_Z_p_O_FDCE ;
input p_desc407_p_O_FDCE ;
input p_ZFF_Y2_8_rep1_Z_p_O_FDCE ;
input p_desc408_p_O_FDCE ;
input p_desc409_p_O_FDCE ;
input p_ZFF_Y2_6_rep1_Z_p_O_FDCE ;
input p_desc410_p_O_FDCE ;
input p_ZFF_Y2_7_rep1_Z_p_O_FDCE ;
input p_desc411_p_O_FDCE ;
input p_ZFF_Y2_14_rep1_Z_p_O_FDCE ;
// instances
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT1 un7_0_10_cry_11_RNO(.I0(ZFF_X1[4:4]),.O(N_2197_i));
defparam un7_0_10_cry_11_RNO.INIT=2'h1;
  LUT1 Y_out_double_2_6_0_cry_0_RNO(.I0(pgZFF_Y1[0:0]),.O(pgZFF_Y1_i));
defparam Y_out_double_2_6_0_cry_0_RNO.INIT=2'h1;
  LUT1 un7_0_6_cry_3_RNO(.I0(ZFF_X1_fast[6:6]),.O(N_3313_i));
defparam un7_0_6_cry_3_RNO.INIT=2'h1;
  LUT1 un6_0_8_cry_21_RNO(.I0(ZFF_X0[11:11]),.O(N_2366_i));
defparam un6_0_8_cry_21_RNO.INIT=2'h1;
  LUT1 desc0(.I0(un9_11_fast[23:23]),.O(un9_11_i[23:23]));
defparam desc0.INIT=2'h1;
  LUT1 un10_8_cry_10_RNO(.I0(ZFF_Y2[5:5]),.O(N_2973_i));
defparam un10_8_cry_10_RNO.INIT=2'h1;
  LUT1 un8_0_8_cry_21_RNO(.I0(ZFF_X2[11:11]),.O(N_3180_i));
defparam un8_0_8_cry_21_RNO.INIT=2'h1;
  LUT1 un6_0_6_cry_3_RNO(.I0(ZFF_X0[8:8]),.O(N_2372_i));
defparam un6_0_6_cry_3_RNO.INIT=2'h1;
  LUT1 un6_0_6_cry_0_RNO(.I0(ZFF_X0[5:5]),.O(N_2379_i));
defparam un6_0_6_cry_0_RNO.INIT=2'h1;
  LUT1 un8_0_6_cry_3_RNO(.I0(ZFF_X2[8:8]),.O(N_3186_i));
defparam un8_0_6_cry_3_RNO.INIT=2'h1;
  LUT1 un8_0_6_cry_0_RNO(.I0(ZFF_X2[5:5]),.O(N_3193_i));
defparam un8_0_6_cry_0_RNO.INIT=2'h1;
  LUT1 un7_0_10_s_27_true_cZ(.I0(GND),.O(un7_0_10_s_27_true));
defparam un7_0_10_s_27_true_cZ.INIT=2'h3;
  LUT2 un9_8_s_36(.I0(un9_8_axb_36),.I1(un9_8[45:45]),.O(un9_8[44:44]));
defparam un9_8_s_36.INIT=4'h6;
  LUT2 un6_0_8_s_27(.I0(un6_0_8_axb_27),.I1(un6_0_8[38:38]),.O(un6_0_8[37:37]));
defparam un6_0_8_s_27.INIT=4'h6;
  LUT2 un8_0_8_s_27(.I0(un8_0_8_axb_27),.I1(un8_0_8[38:38]),.O(un8_0_8[37:37]));
defparam un8_0_8_s_27.INIT=4'h6;
  LUT1 un8_0_8_axb_27_cZ(.I0(GND),.O(un8_0_8_axb_27));
defparam un8_0_8_axb_27_cZ.INIT=2'h3;
  LUT1 un6_0_8_axb_27_cZ(.I0(GND),.O(un6_0_8_axb_27));
defparam un6_0_8_axb_27_cZ.INIT=2'h3;
  LUT1 un9_8_axb_36_cZ(.I0(GND),.O(un9_8_axb_36));
defparam un9_8_axb_36_cZ.INIT=2'h3;
  LUT1 un9_8_axb_35_cZ(.I0(GND),.O(un9_8_axb_35));
defparam un9_8_axb_35_cZ.INIT=2'h3;
  LUT1 un9_8_axb_34_cZ(.I0(GND),.O(un9_8_axb_34));
defparam un9_8_axb_34_cZ.INIT=2'h3;
  LUT1 un9_8_axb_33_cZ(.I0(GND),.O(un9_8_axb_33));
defparam un9_8_axb_33_cZ.INIT=2'h3;
  LUT1 un9_8_axb_32_cZ(.I0(GND),.O(un9_8_axb_32));
defparam un9_8_axb_32_cZ.INIT=2'h3;
  LUT1 un9_8_axb_31_cZ(.I0(GND),.O(un9_8_axb_31));
defparam un9_8_axb_31_cZ.INIT=2'h3;
  LUT1 un7_0_10_axb_26_cZ(.I0(GND),.O(un7_0_10_axb_26));
defparam un7_0_10_axb_26_cZ.INIT=2'h3;
  LD desc1(.Q(pgZFF_Y2_quad[45:45]),.D(un10_s_39),.G(state_reg_ret_5_cb));
defparam desc1.INIT=1'b0;
  LD desc2(.Q(pgZFF_Y2_quad[46:46]),.D(un10_s_40),.G(state_reg_ret_5_cb));
defparam desc2.INIT=1'b0;
  LD desc3(.Q(pgZFF_Y2_quad[47:47]),.D(un10_s_41),.G(state_reg_ret_5_cb));
defparam desc3.INIT=1'b0;
  LD desc4(.Q(pgZFF_Y2_quad[37:37]),.D(un10_s_31),.G(state_reg_ret_5_cb));
defparam desc4.INIT=1'b0;
  LD desc5(.Q(pgZFF_Y2_quad[38:38]),.D(un10_s_32),.G(state_reg_ret_5_cb));
defparam desc5.INIT=1'b0;
  LD desc6(.Q(pgZFF_Y2_quad[39:39]),.D(un10_s_33),.G(state_reg_ret_5_cb));
defparam desc6.INIT=1'b0;
  LD desc7(.Q(pgZFF_Y2_quad[40:40]),.D(un10_s_34),.G(state_reg_ret_5_cb));
defparam desc7.INIT=1'b0;
  LD desc8(.Q(pgZFF_Y2_quad[41:41]),.D(un10_s_35),.G(state_reg_ret_5_cb));
defparam desc8.INIT=1'b0;
  LD desc9(.Q(pgZFF_Y2_quad[42:42]),.D(un10_s_36),.G(state_reg_ret_5_cb));
defparam desc9.INIT=1'b0;
  LD desc10(.Q(pgZFF_Y2_quad[43:43]),.D(un10_s_37),.G(state_reg_ret_5_cb));
defparam desc10.INIT=1'b0;
  LD desc11(.Q(pgZFF_Y2_quad[44:44]),.D(un10_s_38),.G(state_reg_ret_5_cb));
defparam desc11.INIT=1'b0;
  LD desc12(.Q(pgZFF_Y2_quad[30:30]),.D(un10_s_24),.G(state_reg_ret_5_cb));
defparam desc12.INIT=1'b0;
  LD desc13(.Q(pgZFF_Y2_quad[31:31]),.D(un10_s_25),.G(state_reg_ret_5_cb));
defparam desc13.INIT=1'b0;
  LD desc14(.Q(pgZFF_Y2_quad[32:32]),.D(un10_s_26),.G(state_reg_ret_5_cb));
defparam desc14.INIT=1'b0;
  LD desc15(.Q(pgZFF_Y2_quad[33:33]),.D(un10_s_27),.G(state_reg_ret_5_cb));
defparam desc15.INIT=1'b0;
  LD desc16(.Q(pgZFF_Y2_quad[34:34]),.D(un10_s_28),.G(state_reg_ret_5_cb));
defparam desc16.INIT=1'b0;
  LD desc17(.Q(pgZFF_Y2_quad[35:35]),.D(un10_s_29),.G(state_reg_ret_5_cb));
defparam desc17.INIT=1'b0;
  LD desc18(.Q(pgZFF_Y2_quad[36:36]),.D(un10_s_30),.G(state_reg_ret_5_cb));
defparam desc18.INIT=1'b0;
  LD desc19(.Q(pgZFF_Y1_quad[40:40]),.D(un9_s_38),.G(state_reg_ret_5_cb));
defparam desc19.INIT=1'b0;
  LD desc20(.Q(pgZFF_Y1_quad[41:41]),.D(un9_s_39),.G(state_reg_ret_5_cb));
defparam desc20.INIT=1'b0;
  LD desc21(.Q(pgZFF_Y1_quad[42:42]),.D(un9_s_40),.G(state_reg_ret_5_cb));
defparam desc21.INIT=1'b0;
  LD desc22(.Q(pgZFF_Y1_quad[43:43]),.D(un9_s_41),.G(state_reg_ret_5_cb));
defparam desc22.INIT=1'b0;
  LD desc23(.Q(pgZFF_Y1_quad[44:44]),.D(un9_s_42),.G(state_reg_ret_5_cb));
defparam desc23.INIT=1'b0;
  LD desc24(.Q(pgZFF_Y1_quad[45:45]),.D(un9_s_43),.G(state_reg_ret_5_cb));
defparam desc24.INIT=1'b0;
  LD desc25(.Q(pgZFF_Y1_quad[46:46]),.D(un9_s_44),.G(state_reg_ret_5_cb));
defparam desc25.INIT=1'b0;
  LD desc26(.Q(pgZFF_Y1_quad[47:47]),.D(un9_s_45),.G(state_reg_ret_5_cb));
defparam desc26.INIT=1'b0;
  LD desc27(.Q(pgZFF_Y1_quad[33:33]),.D(un9_s_31),.G(state_reg_ret_5_cb));
defparam desc27.INIT=1'b0;
  LD desc28(.Q(pgZFF_Y1_quad[34:34]),.D(un9_s_32),.G(state_reg_ret_5_cb));
defparam desc28.INIT=1'b0;
  LD desc29(.Q(pgZFF_Y1_quad[35:35]),.D(un9_s_33),.G(state_reg_ret_5_cb));
defparam desc29.INIT=1'b0;
  LD desc30(.Q(pgZFF_Y1_quad[36:36]),.D(un9_s_34),.G(state_reg_ret_5_cb));
defparam desc30.INIT=1'b0;
  LD desc31(.Q(pgZFF_Y1_quad[37:37]),.D(un9_s_35),.G(state_reg_ret_5_cb));
defparam desc31.INIT=1'b0;
  LD desc32(.Q(pgZFF_Y1_quad[38:38]),.D(un9_s_36),.G(state_reg_ret_5_cb));
defparam desc32.INIT=1'b0;
  LD desc33(.Q(pgZFF_Y1_quad[39:39]),.D(un9_s_37),.G(state_reg_ret_5_cb));
defparam desc33.INIT=1'b0;
  LD desc34(.Q(pgZFF_X2_quad[42:42]),.D(un8_0_0_s_40),.G(state_reg_ret_5_cb));
defparam desc34.INIT=1'b0;
  LD desc35(.Q(pgZFF_X2_quad[43:43]),.D(un8_0_0_s_41),.G(state_reg_ret_5_cb));
defparam desc35.INIT=1'b0;
  LD desc36(.Q(pgZFF_X2_quad[44:44]),.D(un8_0_0_s_42),.G(state_reg_ret_5_cb));
defparam desc36.INIT=1'b0;
  LD desc37(.Q(pgZFF_X2_quad[46:46]),.D(un8_0_0_s_43),.G(state_reg_ret_5_cb));
defparam desc37.INIT=1'b0;
  LD desc38(.Q(pgZFF_Y1_quad[30:30]),.D(un9_s_28),.G(state_reg_ret_5_cb));
defparam desc38.INIT=1'b0;
  LD desc39(.Q(pgZFF_Y1_quad[31:31]),.D(un9_s_29),.G(state_reg_ret_5_cb));
defparam desc39.INIT=1'b0;
  LD desc40(.Q(pgZFF_Y1_quad[32:32]),.D(un9_s_30),.G(state_reg_ret_5_cb));
defparam desc40.INIT=1'b0;
  LD desc41(.Q(pgZFF_X2_quad[35:35]),.D(un8_0_0_s_33),.G(state_reg_ret_5_cb));
defparam desc41.INIT=1'b0;
  LD desc42(.Q(pgZFF_X2_quad[36:36]),.D(un8_0_0_s_34),.G(state_reg_ret_5_cb));
defparam desc42.INIT=1'b0;
  LD desc43(.Q(pgZFF_X2_quad[37:37]),.D(un8_0_0_s_35),.G(state_reg_ret_5_cb));
defparam desc43.INIT=1'b0;
  LD desc44(.Q(pgZFF_X2_quad[38:38]),.D(un8_0_0_s_36),.G(state_reg_ret_5_cb));
defparam desc44.INIT=1'b0;
  LD desc45(.Q(pgZFF_X2_quad[39:39]),.D(un8_0_0_s_37),.G(state_reg_ret_5_cb));
defparam desc45.INIT=1'b0;
  LD desc46(.Q(pgZFF_X2_quad[40:40]),.D(un8_0_0_s_38),.G(state_reg_ret_5_cb));
defparam desc46.INIT=1'b0;
  LD desc47(.Q(pgZFF_X2_quad[41:41]),.D(un8_0_0_s_39),.G(state_reg_ret_5_cb));
defparam desc47.INIT=1'b0;
  LD desc48(.Q(pgZFF_X1_quad[45:45]),.D(un7_0_0_s_44),.G(state_reg_ret_5_cb));
defparam desc48.INIT=1'b0;
  LD desc49(.Q(pgZFF_X1_quad[47:47]),.D(un7_0_0_s_45),.G(state_reg_ret_5_cb));
defparam desc49.INIT=1'b0;
  LD desc50(.Q(pgZFF_X2_quad[30:30]),.D(un8_0_0_s_28),.G(state_reg_ret_5_cb));
defparam desc50.INIT=1'b0;
  LD desc51(.Q(pgZFF_X2_quad[31:31]),.D(un8_0_0_s_29),.G(state_reg_ret_5_cb));
defparam desc51.INIT=1'b0;
  LD desc52(.Q(pgZFF_X2_quad[32:32]),.D(un8_0_0_s_30),.G(state_reg_ret_5_cb));
defparam desc52.INIT=1'b0;
  LD desc53(.Q(pgZFF_X2_quad[33:33]),.D(un8_0_0_s_31),.G(state_reg_ret_5_cb));
defparam desc53.INIT=1'b0;
  LD desc54(.Q(pgZFF_X2_quad[34:34]),.D(un8_0_0_s_32),.G(state_reg_ret_5_cb));
defparam desc54.INIT=1'b0;
  LD desc55(.Q(pgZFF_X1_quad[38:38]),.D(un7_0_0_s_37),.G(state_reg_ret_5_cb));
defparam desc55.INIT=1'b0;
  LD desc56(.Q(pgZFF_X1_quad[39:39]),.D(un7_0_0_s_38),.G(state_reg_ret_5_cb));
defparam desc56.INIT=1'b0;
  LD desc57(.Q(pgZFF_X1_quad[40:40]),.D(un7_0_0_s_39),.G(state_reg_ret_5_cb));
defparam desc57.INIT=1'b0;
  LD desc58(.Q(pgZFF_X1_quad[41:41]),.D(un7_0_0_s_40),.G(state_reg_ret_5_cb));
defparam desc58.INIT=1'b0;
  LD desc59(.Q(pgZFF_X1_quad[42:42]),.D(un7_0_0_s_41),.G(state_reg_ret_5_cb));
defparam desc59.INIT=1'b0;
  LD desc60(.Q(pgZFF_X1_quad[43:43]),.D(un7_0_0_s_42),.G(state_reg_ret_5_cb));
defparam desc60.INIT=1'b0;
  LD desc61(.Q(pgZFF_X1_quad[44:44]),.D(un7_0_0_s_43),.G(state_reg_ret_5_cb));
defparam desc61.INIT=1'b0;
  LD desc62(.Q(pgZFF_X1_quad[30:30]),.D(un7_0_0_s_29),.G(state_reg_ret_5_cb));
defparam desc62.INIT=1'b0;
  LD desc63(.Q(pgZFF_X1_quad[31:31]),.D(un7_0_0_s_30),.G(state_reg_ret_5_cb));
defparam desc63.INIT=1'b0;
  LD desc64(.Q(pgZFF_X1_quad[32:32]),.D(un7_0_0_s_31),.G(state_reg_ret_5_cb));
defparam desc64.INIT=1'b0;
  LD desc65(.Q(pgZFF_X1_quad[33:33]),.D(un7_0_0_s_32),.G(state_reg_ret_5_cb));
defparam desc65.INIT=1'b0;
  LD desc66(.Q(pgZFF_X1_quad[34:34]),.D(un7_0_0_s_33),.G(state_reg_ret_5_cb));
defparam desc66.INIT=1'b0;
  LD desc67(.Q(pgZFF_X1_quad[35:35]),.D(un7_0_0_s_34),.G(state_reg_ret_5_cb));
defparam desc67.INIT=1'b0;
  LD desc68(.Q(pgZFF_X1_quad[36:36]),.D(un7_0_0_s_35),.G(state_reg_ret_5_cb));
defparam desc68.INIT=1'b0;
  LD desc69(.Q(pgZFF_X1_quad[37:37]),.D(un7_0_0_s_36),.G(state_reg_ret_5_cb));
defparam desc69.INIT=1'b0;
  LD desc70(.Q(pgZFF_X0_quad[40:40]),.D(un6_0_0_s_38),.G(state_reg_ret_5_cb));
defparam desc70.INIT=1'b0;
  LD desc71(.Q(pgZFF_X0_quad[41:41]),.D(un6_0_0_s_39),.G(state_reg_ret_5_cb));
defparam desc71.INIT=1'b0;
  LD desc72(.Q(pgZFF_X0_quad[42:42]),.D(un6_0_0_s_40),.G(state_reg_ret_5_cb));
defparam desc72.INIT=1'b0;
  LD desc73(.Q(pgZFF_X0_quad[43:43]),.D(un6_0_0_s_41),.G(state_reg_ret_5_cb));
defparam desc73.INIT=1'b0;
  LD desc74(.Q(pgZFF_X0_quad[44:44]),.D(un6_0_0_s_42),.G(state_reg_ret_5_cb));
defparam desc74.INIT=1'b0;
  LD desc75(.Q(pgZFF_X0_quad[46:46]),.D(un6_0_0_s_43),.G(state_reg_ret_5_cb));
defparam desc75.INIT=1'b0;
  LD desc76(.Q(pgZFF_X0_quad[32:32]),.D(un6_0_0_s_30),.G(state_reg_ret_5_cb));
defparam desc76.INIT=1'b0;
  LD desc77(.Q(pgZFF_X0_quad[33:33]),.D(un6_0_0_s_31),.G(state_reg_ret_5_cb));
defparam desc77.INIT=1'b0;
  LD desc78(.Q(pgZFF_X0_quad[34:34]),.D(un6_0_0_s_32),.G(state_reg_ret_5_cb));
defparam desc78.INIT=1'b0;
  LD desc79(.Q(pgZFF_X0_quad[35:35]),.D(un6_0_0_s_33),.G(state_reg_ret_5_cb));
defparam desc79.INIT=1'b0;
  LD desc80(.Q(pgZFF_X0_quad[36:36]),.D(un6_0_0_s_34),.G(state_reg_ret_5_cb));
defparam desc80.INIT=1'b0;
  LD desc81(.Q(pgZFF_X0_quad[37:37]),.D(un6_0_0_s_35),.G(state_reg_ret_5_cb));
defparam desc81.INIT=1'b0;
  LD desc82(.Q(pgZFF_X0_quad[38:38]),.D(un6_0_0_s_36),.G(state_reg_ret_5_cb));
defparam desc82.INIT=1'b0;
  LD desc83(.Q(pgZFF_X0_quad[39:39]),.D(un6_0_0_s_37),.G(state_reg_ret_5_cb));
defparam desc83.INIT=1'b0;
  LD desc84(.Q(pgZFF_X0_quad[30:30]),.D(un6_0_0_s_28),.G(state_reg_ret_5_cb));
defparam desc84.INIT=1'b0;
  LD desc85(.Q(pgZFF_X0_quad[31:31]),.D(un6_0_0_s_29),.G(state_reg_ret_5_cb));
defparam desc85.INIT=1'b0;
  p_O_FDE desc86(.Q(pgZFF_Y1[17:17]),.D(pgZFF_Y1_quad[47:47]),.C(clk),.CE(trunc_prods),.E(p_desc86_p_O_FDE));
defparam desc86.INIT=1'b0;
  p_O_FDE desc87(.Q(pgZFF_Y1[16:16]),.D(pgZFF_Y1_quad[46:46]),.C(clk),.CE(trunc_prods),.E(p_desc87_p_O_FDE));
defparam desc87.INIT=1'b0;
  p_O_FDE desc88(.Q(pgZFF_Y1[15:15]),.D(pgZFF_Y1_quad[45:45]),.C(clk),.CE(trunc_prods),.E(p_desc88_p_O_FDE));
defparam desc88.INIT=1'b0;
  p_O_FDE desc89(.Q(pgZFF_Y1[14:14]),.D(pgZFF_Y1_quad[44:44]),.C(clk),.CE(trunc_prods),.E(p_desc89_p_O_FDE));
defparam desc89.INIT=1'b0;
  p_O_FDE desc90(.Q(pgZFF_Y1[13:13]),.D(pgZFF_Y1_quad[43:43]),.C(clk),.CE(trunc_prods),.E(p_desc90_p_O_FDE));
defparam desc90.INIT=1'b0;
  p_O_FDE desc91(.Q(pgZFF_Y1[12:12]),.D(pgZFF_Y1_quad[42:42]),.C(clk),.CE(trunc_prods),.E(p_desc91_p_O_FDE));
defparam desc91.INIT=1'b0;
  p_O_FDE desc92(.Q(pgZFF_Y1[11:11]),.D(pgZFF_Y1_quad[41:41]),.C(clk),.CE(trunc_prods),.E(p_desc92_p_O_FDE));
defparam desc92.INIT=1'b0;
  p_O_FDE desc93(.Q(pgZFF_Y1[10:10]),.D(pgZFF_Y1_quad[40:40]),.C(clk),.CE(trunc_prods),.E(p_desc93_p_O_FDE));
defparam desc93.INIT=1'b0;
  p_O_FDE desc94(.Q(pgZFF_Y1[9:9]),.D(pgZFF_Y1_quad[39:39]),.C(clk),.CE(trunc_prods),.E(p_desc94_p_O_FDE));
defparam desc94.INIT=1'b0;
  p_O_FDE desc95(.Q(pgZFF_Y1[8:8]),.D(pgZFF_Y1_quad[38:38]),.C(clk),.CE(trunc_prods),.E(p_desc95_p_O_FDE));
defparam desc95.INIT=1'b0;
  p_O_FDE desc96(.Q(pgZFF_Y1[7:7]),.D(pgZFF_Y1_quad[37:37]),.C(clk),.CE(trunc_prods),.E(p_desc96_p_O_FDE));
defparam desc96.INIT=1'b0;
  p_O_FDE desc97(.Q(pgZFF_Y1[6:6]),.D(pgZFF_Y1_quad[36:36]),.C(clk),.CE(trunc_prods),.E(p_desc97_p_O_FDE));
defparam desc97.INIT=1'b0;
  p_O_FDE desc98(.Q(pgZFF_Y1[5:5]),.D(pgZFF_Y1_quad[35:35]),.C(clk),.CE(trunc_prods),.E(p_desc98_p_O_FDE));
defparam desc98.INIT=1'b0;
  p_O_FDE desc99(.Q(pgZFF_Y1[4:4]),.D(pgZFF_Y1_quad[34:34]),.C(clk),.CE(trunc_prods),.E(p_desc99_p_O_FDE));
defparam desc99.INIT=1'b0;
  p_O_FDE desc100(.Q(pgZFF_Y1[3:3]),.D(pgZFF_Y1_quad[33:33]),.C(clk),.CE(trunc_prods),.E(p_desc100_p_O_FDE));
defparam desc100.INIT=1'b0;
  p_O_FDE desc101(.Q(pgZFF_Y1[2:2]),.D(pgZFF_Y1_quad[32:32]),.C(clk),.CE(trunc_prods),.E(p_desc101_p_O_FDE));
defparam desc101.INIT=1'b0;
  p_O_FDE desc102(.Q(pgZFF_Y1[1:1]),.D(pgZFF_Y1_quad[31:31]),.C(clk),.CE(trunc_prods),.E(p_desc102_p_O_FDE));
defparam desc102.INIT=1'b0;
  p_O_FDE desc103(.Q(pgZFF_Y1[0:0]),.D(pgZFF_Y1_quad[30:30]),.C(clk),.CE(trunc_prods),.E(p_desc103_p_O_FDE));
defparam desc103.INIT=1'b0;
  p_O_FDE desc104(.Q(pgZFF_Y2[17:17]),.D(pgZFF_Y2_quad[47:47]),.C(clk),.CE(trunc_prods),.E(p_desc104_p_O_FDE));
defparam desc104.INIT=1'b0;
  p_O_FDE desc105(.Q(pgZFF_Y2[16:16]),.D(pgZFF_Y2_quad[46:46]),.C(clk),.CE(trunc_prods),.E(p_desc105_p_O_FDE));
defparam desc105.INIT=1'b0;
  p_O_FDE desc106(.Q(pgZFF_Y2[15:15]),.D(pgZFF_Y2_quad[45:45]),.C(clk),.CE(trunc_prods),.E(p_desc106_p_O_FDE));
defparam desc106.INIT=1'b0;
  p_O_FDE desc107(.Q(pgZFF_Y2[14:14]),.D(pgZFF_Y2_quad[44:44]),.C(clk),.CE(trunc_prods),.E(p_desc107_p_O_FDE));
defparam desc107.INIT=1'b0;
  p_O_FDE desc108(.Q(pgZFF_Y2[13:13]),.D(pgZFF_Y2_quad[43:43]),.C(clk),.CE(trunc_prods),.E(p_desc108_p_O_FDE));
defparam desc108.INIT=1'b0;
  p_O_FDE desc109(.Q(pgZFF_Y2[12:12]),.D(pgZFF_Y2_quad[42:42]),.C(clk),.CE(trunc_prods),.E(p_desc109_p_O_FDE));
defparam desc109.INIT=1'b0;
  p_O_FDE desc110(.Q(pgZFF_Y2[11:11]),.D(pgZFF_Y2_quad[41:41]),.C(clk),.CE(trunc_prods),.E(p_desc110_p_O_FDE));
defparam desc110.INIT=1'b0;
  p_O_FDE desc111(.Q(pgZFF_Y2[10:10]),.D(pgZFF_Y2_quad[40:40]),.C(clk),.CE(trunc_prods),.E(p_desc111_p_O_FDE));
defparam desc111.INIT=1'b0;
  p_O_FDE desc112(.Q(pgZFF_Y2[9:9]),.D(pgZFF_Y2_quad[39:39]),.C(clk),.CE(trunc_prods),.E(p_desc112_p_O_FDE));
defparam desc112.INIT=1'b0;
  p_O_FDE desc113(.Q(pgZFF_Y2[8:8]),.D(pgZFF_Y2_quad[38:38]),.C(clk),.CE(trunc_prods),.E(p_desc113_p_O_FDE));
defparam desc113.INIT=1'b0;
  p_O_FDE desc114(.Q(pgZFF_Y2[7:7]),.D(pgZFF_Y2_quad[37:37]),.C(clk),.CE(trunc_prods),.E(p_desc114_p_O_FDE));
defparam desc114.INIT=1'b0;
  p_O_FDE desc115(.Q(pgZFF_Y2[6:6]),.D(pgZFF_Y2_quad[36:36]),.C(clk),.CE(trunc_prods),.E(p_desc115_p_O_FDE));
defparam desc115.INIT=1'b0;
  p_O_FDE desc116(.Q(pgZFF_Y2[5:5]),.D(pgZFF_Y2_quad[35:35]),.C(clk),.CE(trunc_prods),.E(p_desc116_p_O_FDE));
defparam desc116.INIT=1'b0;
  p_O_FDE desc117(.Q(pgZFF_Y2[4:4]),.D(pgZFF_Y2_quad[34:34]),.C(clk),.CE(trunc_prods),.E(p_desc117_p_O_FDE));
defparam desc117.INIT=1'b0;
  p_O_FDE desc118(.Q(pgZFF_Y2[3:3]),.D(pgZFF_Y2_quad[33:33]),.C(clk),.CE(trunc_prods),.E(p_desc118_p_O_FDE));
defparam desc118.INIT=1'b0;
  p_O_FDE desc119(.Q(pgZFF_Y2[2:2]),.D(pgZFF_Y2_quad[32:32]),.C(clk),.CE(trunc_prods),.E(p_desc119_p_O_FDE));
defparam desc119.INIT=1'b0;
  p_O_FDE desc120(.Q(pgZFF_Y2[1:1]),.D(pgZFF_Y2_quad[31:31]),.C(clk),.CE(trunc_prods),.E(p_desc120_p_O_FDE));
defparam desc120.INIT=1'b0;
  p_O_FDE desc121(.Q(pgZFF_Y2[0:0]),.D(pgZFF_Y2_quad[30:30]),.C(clk),.CE(trunc_prods),.E(p_desc121_p_O_FDE));
defparam desc121.INIT=1'b0;
  LUT3 ZFF_X1_10_rep1_RNIEAHH(.I0(ZFF_X1[9:9]),.I1(ZFF_X1_10_rep1),.I2(ZFF_X1_15_rep1),.O(un7_0_10_axb_1));
defparam ZFF_X1_10_rep1_RNIEAHH.INIT=8'h6C;
  LUT1 un7_0_10_axb_2_cZ(.I0(ZFF_X1_11_rep1),.O(un7_0_10_axb_2));
defparam un7_0_10_axb_2_cZ.INIT=2'h2;
  LUT1 un7_0_10_axb_3_cZ(.I0(ZFF_X1[12:12]),.O(un7_0_10_axb_3));
defparam un7_0_10_axb_3_cZ.INIT=2'h2;
  LUT2 un7_0_10_axb_4_cZ(.I0(ZFF_X1[16:16]),.I1(ZFF_X1_13_rep1),.O(un7_0_10_axb_4));
defparam un7_0_10_axb_4_cZ.INIT=4'h6;
  LUT2 un7_0_10_axb_5_cZ(.I0(ZFF_X1[14:14]),.I1(ZFF_X1[16:16]),.O(un7_0_10_axb_5));
defparam un7_0_10_axb_5_cZ.INIT=4'h6;
  LUT2 un7_0_10_axb_6_cZ(.I0(ZFF_X1[15:15]),.I1(ZFF_X1[16:16]),.O(un7_0_10_axb_6));
defparam un7_0_10_axb_6_cZ.INIT=4'h6;
  LUT1 un7_0_10_axb_7_cZ(.I0(ZFF_X1[0:0]),.O(un7_0_10_axb_7));
defparam un7_0_10_axb_7_cZ.INIT=2'h1;
  LUT1 un7_0_10_axb_8_cZ(.I0(ZFF_X1[1:1]),.O(un7_0_10_axb_8));
defparam un7_0_10_axb_8_cZ.INIT=2'h1;
  LUT1 un7_0_10_axb_9_cZ(.I0(ZFF_X1[2:2]),.O(un7_0_10_axb_9));
defparam un7_0_10_axb_9_cZ.INIT=2'h1;
  LUT2 un7_0_10_axb_10_cZ(.I0(ZFF_X1[0:0]),.I1(ZFF_X1[3:3]),.O(un7_0_10_axb_10));
defparam un7_0_10_axb_10_cZ.INIT=4'h9;
  LUT3 un7_0_10_axb_11_cZ(.I0(ZFF_X1[1:1]),.I1(ZFF_X1[4:4]),.I2(ZFF_X1[16:16]),.O(un7_0_10_axb_11));
defparam un7_0_10_axb_11_cZ.INIT=8'h69;
  LUT4 desc122(.I0(ZFF_X1[1:1]),.I1(ZFF_X1[2:2]),.I2(ZFF_X1[5:5]),.I3(ZFF_X1[16:16]),.O(un7_0_10_axb_12));
defparam desc122.INIT=16'h69C3;
  LUT4 un7_0_10_axb_16_cZ(.I0(ZFF_X1[5:5]),.I1(ZFF_X1[6:6]),.I2(ZFF_X1[8:8]),.I3(ZFF_X1[9:9]),.O(un7_0_10_axb_16));
defparam un7_0_10_axb_16_cZ.INIT=16'h9C63;
  LUT4 un7_0_10_axb_17_cZ(.I0(ZFF_X1[6:6]),.I1(ZFF_X1[7:7]),.I2(ZFF_X1[9:9]),.I3(ZFF_X1[10:10]),.O(un7_0_10_axb_17));
defparam un7_0_10_axb_17_cZ.INIT=16'h9C63;
  LUT4 un7_0_10_axb_18_cZ(.I0(ZFF_X1[7:7]),.I1(ZFF_X1[8:8]),.I2(ZFF_X1[10:10]),.I3(ZFF_X1[11:11]),.O(un7_0_10_axb_18));
defparam un7_0_10_axb_18_cZ.INIT=16'h9C63;
  LUT4 un7_0_10_axb_19_cZ(.I0(ZFF_X1[8:8]),.I1(ZFF_X1[9:9]),.I2(ZFF_X1[11:11]),.I3(ZFF_X1[12:12]),.O(un7_0_10_axb_19));
defparam un7_0_10_axb_19_cZ.INIT=16'h9C63;
  LUT4 un7_0_10_axb_20_cZ(.I0(ZFF_X1[9:9]),.I1(ZFF_X1[10:10]),.I2(ZFF_X1[12:12]),.I3(ZFF_X1[13:13]),.O(un7_0_10_axb_20));
defparam un7_0_10_axb_20_cZ.INIT=16'h9C63;
  LUT4 un7_0_10_axb_21_cZ(.I0(ZFF_X1[10:10]),.I1(ZFF_X1[11:11]),.I2(ZFF_X1[13:13]),.I3(ZFF_X1[14:14]),.O(un7_0_10_axb_21));
defparam un7_0_10_axb_21_cZ.INIT=16'h9C63;
  LUT4 un7_0_10_axb_22_cZ(.I0(ZFF_X1[11:11]),.I1(ZFF_X1[12:12]),.I2(ZFF_X1[14:14]),.I3(ZFF_X1[15:15]),.O(un7_0_10_axb_22));
defparam un7_0_10_axb_22_cZ.INIT=16'h9C63;
  LUT3 un7_0_10_axb_23_cZ(.I0(ZFF_X1[12:12]),.I1(ZFF_X1[13:13]),.I2(ZFF_X1[15:15]),.O(un7_0_10_axb_23));
defparam un7_0_10_axb_23_cZ.INIT=8'h63;
  LUT1 desc123(.I0(ZFF_X1[14:14]),.O(N_3387_i));
defparam desc123.INIT=2'h1;
  LUT1 desc124(.I0(ZFF_X1[15:15]),.O(N_3385_i));
defparam desc124.INIT=2'h1;
  LUT1 un6_0_0_cry_0_RNO(.I0(ZFF_X0[0:0]),.O(N_2393_i));
defparam un6_0_0_cry_0_RNO.INIT=2'h1;
  LUT1 un6_0_0_cry_1_RNO(.I0(ZFF_X0[1:1]),.O(N_2390_i));
defparam un6_0_0_cry_1_RNO.INIT=2'h1;
  LUT1 un6_0_0_cry_2_RNO(.I0(ZFF_X0[2:2]),.O(N_2387_i));
defparam un6_0_0_cry_2_RNO.INIT=2'h1;
  LUT1 un6_0_0_cry_3_RNO(.I0(ZFF_X0[3:3]),.O(N_2384_i));
defparam un6_0_0_cry_3_RNO.INIT=2'h1;
  LUT1 un6_0_0_cry_4_RNO(.I0(ZFF_X0[4:4]),.O(N_2381_i));
defparam un6_0_0_cry_4_RNO.INIT=2'h1;
  LUT2 un6_0_0_cry_5_RNO(.I0(ZFF_X0[0:0]),.I1(ZFF_X0[5:5]),.O(un6_0_6[5:5]));
defparam un6_0_0_cry_5_RNO.INIT=4'h9;
  LUT1 un6_0_0_cry_6_RNO(.I0(un6_0_6[6:6]),.O(un6_0_0_cry_6_sf));
defparam un6_0_0_cry_6_RNO.INIT=2'h2;
  LUT2 un6_0_0_axb_7_cZ(.I0(ZFF_X0[2:2]),.I1(un6_0_6[7:7]),.O(un6_0_0_axb_7));
defparam un6_0_0_axb_7_cZ.INIT=4'h6;
  LUT2 un6_0_0_axb_8_cZ(.I0(ZFF_X0[0:0]),.I1(un6_0_6[8:8]),.O(un6_0_0_axb_8));
defparam un6_0_0_axb_8_cZ.INIT=4'h6;
  LUT2 un6_0_0_axb_9_cZ(.I0(ZFF_X0[1:1]),.I1(un6_0_6[9:9]),.O(un6_0_0_axb_9));
defparam un6_0_0_axb_9_cZ.INIT=4'h6;
  LUT3 un6_0_0_axb_10_cZ(.I0(ZFF_X0[2:2]),.I1(ZFF_X0[3:3]),.I2(un6_0_6[10:10]),.O(un6_0_0_axb_10));
defparam un6_0_0_axb_10_cZ.INIT=8'h96;
  LUT4 un6_0_0_axb_12_cZ(.I0(un6_0_6[11:11]),.I1(un6_0_6[12:12]),.I2(un6_0_8[11:11]),.I3(un6_0_8[12:12]),.O(un6_0_0_axb_12));
defparam un6_0_0_axb_12_cZ.INIT=16'h936C;
  LUT4 un6_0_0_axb_13_cZ(.I0(un6_0_6[12:12]),.I1(un6_0_6[13:13]),.I2(un6_0_8[12:12]),.I3(un6_0_8[13:13]),.O(un6_0_0_axb_13));
defparam un6_0_0_axb_13_cZ.INIT=16'h936C;
  LUT4 un6_0_0_axb_14_cZ(.I0(un6_0_6[13:13]),.I1(un6_0_6[14:14]),.I2(un6_0_8[13:13]),.I3(un6_0_8[14:14]),.O(un6_0_0_axb_14));
defparam un6_0_0_axb_14_cZ.INIT=16'h936C;
  LUT4 un6_0_9_s_15_RNIP1BU(.I0(un6_0_8[29:29]),.I1(un6_0_8[30:30]),.I2(un6_0_9[29:29]),.I3(un6_0_9[30:30]),.O(un6_0_0_axb_30));
defparam un6_0_9_s_15_RNIP1BU.INIT=16'h936C;
  LUT4 un6_0_9_s_15_RNIK2BU(.I0(un6_0_8[30:30]),.I1(un6_0_8[31:31]),.I2(un6_0_9[30:30]),.I3(un6_0_9[31:31]),.O(un6_0_0_axb_31));
defparam un6_0_9_s_15_RNIK2BU.INIT=16'h936C;
  LUT4 un6_0_9_s_16_RNIO2BU(.I0(un6_0_8[31:31]),.I1(un6_0_8[32:32]),.I2(un6_0_9[31:31]),.I3(un6_0_9[32:32]),.O(un6_0_0_axb_32));
defparam un6_0_9_s_16_RNIO2BU.INIT=16'h936C;
  LUT4 un6_0_9_s_17_RNIS2BU(.I0(un6_0_8[32:32]),.I1(un6_0_8[33:33]),.I2(un6_0_9[32:32]),.I3(un6_0_9[33:33]),.O(un6_0_0_axb_33));
defparam un6_0_9_s_17_RNIS2BU.INIT=16'h936C;
  LUT4 un6_0_9_s_18_RNI03BU(.I0(un6_0_8[33:33]),.I1(un6_0_8[34:34]),.I2(un6_0_9[33:33]),.I3(un6_0_9[34:34]),.O(un6_0_0_axb_34));
defparam un6_0_9_s_18_RNI03BU.INIT=16'h936C;
  LUT4 un6_0_9_s_19_RNIR3BU(.I0(un6_0_8[34:34]),.I1(un6_0_8[35:35]),.I2(un6_0_9[34:34]),.I3(un6_0_9[35:35]),.O(un6_0_0_axb_35));
defparam un6_0_9_s_19_RNIR3BU.INIT=16'h936C;
  LUT2 un6_0_6_cry_0_RNO_0(.I0(ZFF_X0[0:0]),.I1(ZFF_X0[5:5]),.O(un6_0_6_cry_0_sf));
defparam un6_0_6_cry_0_RNO_0.INIT=4'h9;
  LUT2 ZFF_X0_1_rep1_RNIF489(.I0(ZFF_X0[6:6]),.I1(ZFF_X0_1_rep1),.O(un6_0_6_axb_1));
defparam ZFF_X0_1_rep1_RNIF489.INIT=4'h9;
  LUT2 desc125(.I0(ZFF_X0[0:0]),.I1(ZFF_X0[7:7]),.O(un6_0_6_axb_2));
defparam desc125.INIT=4'h9;
  LUT3 un6_0_6_axb_3_cZ(.I0(ZFF_X0[8:8]),.I1(ZFF_X0_1_rep1),.I2(ZFF_X0_3_rep1),.O(un6_0_6_axb_3));
defparam un6_0_6_axb_3_cZ.INIT=8'h69;
  LUT4 ZFF_X0_14_rep1_RNI231I1(.I0(ZFF_X0[12:12]),.I1(ZFF_X0[13:13]),.I2(ZFF_X0_14_rep1),.I3(ZFF_X0_15_rep1),.O(un6_0_6_axb_20));
defparam ZFF_X0_14_rep1_RNI231I1.INIT=16'h936C;
  LUT3 desc126(.I0(ZFF_X0[13:13]),.I1(ZFF_X0[14:14]),.I2(ZFF_X0[15:15]),.O(un6_0_6_axb_21));
defparam desc126.INIT=8'h6C;
  LUT1 un6_0_6_axb_22_cZ(.I0(ZFF_X0[15:15]),.O(un6_0_6_axb_22));
defparam un6_0_6_axb_22_cZ.INIT=2'h2;
  LUT2 desc127(.I0(pgZFF_Y1[0:0]),.I1(pgZFF_Y2[0:0]),.O(Y_out_double_2_6_0_axb_0));
defparam desc127.INIT=4'h6;
  LUT3 Y_out_double_2_6_0_axb_1_cZ(.I0(pgZFF_X1[1:1]),.I1(pgZFF_Y1[1:1]),.I2(pgZFF_Y2[1:1]),.O(Y_out_double_2_6_0_axb_1));
defparam Y_out_double_2_6_0_axb_1_cZ.INIT=8'h96;
  LUT2 un9_6_cZ(.I0(un9_8[7:7]),.I1(un9_10[8:8]),.O(un9_6[2:2]));
defparam un9_6_cZ.INIT=4'h9;
  LUT2 un9_axb_4_cZ(.I0(un9_6[6:6]),.I1(un9_8[6:6]),.O(un9_axb_4));
defparam un9_axb_4_cZ.INIT=4'h6;
  LUT2 un9_axb_5_cZ(.I0(un9_6[7:7]),.I1(un9_8[7:7]),.O(un9_axb_5));
defparam un9_axb_5_cZ.INIT=4'h6;
  LUT4 un9_axb_6_cZ(.I0(ZFF_Y1[3:3]),.I1(ZFF_Y1[6:6]),.I2(un9_6[8:8]),.I3(un9_10[8:8]),.O(un9_axb_6));
defparam un9_axb_6_cZ.INIT=16'h9669;
  LUT4 un9_8_s_36_RNIA8E41(.I0(un9_6[43:43]),.I1(un9_6[44:44]),.I2(un9_8[43:43]),.I3(un9_8[44:44]),.O(un9_axb_42));
defparam un9_8_s_36_RNIA8E41.INIT=16'h936C;
  LUT4 un9_8_s_36_RNI7SF81(.I0(un9_6[44:44]),.I1(un9_6[45:45]),.I2(un9_8[44:44]),.I3(un9_8[45:45]),.O(un9_axb_43));
defparam un9_8_s_36_RNI7SF81.INIT=16'h6C93;
  LUT4 un9_8_cry_37_outext_RNIDUB71(.I0(un9_6[45:45]),.I1(un9_6[46:46]),.I2(un9_8[45:45]),.I3(un9_8[46:46]),.O(un9_axb_44));
defparam un9_8_cry_37_outext_RNIDUB71.INIT=16'h39C6;
  LUT4 desc128(.I0(ZFF_Y1_4_rep1),.I1(ZFF_Y1_5_rep1),.I2(ZFF_Y1_fast[6:6]),.I3(un9_10_8_rep1),.O(un9_6_0_axb_6));
defparam desc128.INIT=16'h695A;
  LUT4 desc129(.I0(ZFF_Y1_4_rep1),.I1(ZFF_Y1_5_rep1),.I2(ZFF_Y1_fast[6:6]),.I3(ZFF_Y1_fast[7:7]),.O(un9_6_0_axb_7));
defparam desc129.INIT=16'h36C9;
  LUT1 un9_6_0_cry_9_RNO_cZ(.I0(ZFF_Y1_9_rep1),.O(un9_6_0_cry_9_RNO));
defparam un9_6_0_cry_9_RNO_cZ.INIT=2'h1;
  LUT2 un9_6_24(.I0(un9_10_8_rep1),.I1(un9_11_22_rep1),.O(un9_6_0_axb_10));
defparam un9_6_24.INIT=4'h9;
  LUT4 ZFF_Y1_10_rep1_RNI7IP21(.I0(un9_8_6_rep1),.I1(un9_10_8_rep1),.I2(un9_11_22_rep1),.I3(un9_11_fast[23:23]),.O(un9_6_0_axb_11));
defparam ZFF_Y1_10_rep1_RNI7IP21.INIT=16'hA659;
  LUT4 ZFF_Y1_1_rep1_RNIDGMG1(.I0(ZFF_Y1_4_rep1),.I1(un9_8_6_rep1),.I2(un9_11_24_rep1),.I3(un9_11_fast[23:23]),.O(un9_6_0_axb_12));
defparam ZFF_Y1_1_rep1_RNIDGMG1.INIT=16'hA569;
  LUT4 desc130(.I0(ZFF_Y1[5:5]),.I1(ZFF_Y1_4_rep1),.I2(un9_11_24_rep1),.I3(un9_11_25_rep1),.O(un9_6_0_axb_13));
defparam desc130.INIT=16'hA659;
  LUT4 ZFF_Y1_14_rep1_RNILL101(.I0(ZFF_Y1_5_rep1),.I1(un9_11_24_rep1),.I2(un9_11_25_rep1),.I3(un9_11_26_rep1),.O(un9_6_0_axb_14));
defparam ZFF_Y1_14_rep1_RNILL101.INIT=16'h39C6;
  LUT4 ZFF_Y1_10_rep1_RNI3S241(.I0(ZFF_Y1_15_rep1),.I1(un9_11_22_rep1),.I2(un9_11_24_rep1),.I3(un9_11_26_rep1),.O(un9_6_0_axb_15));
defparam ZFF_Y1_10_rep1_RNI3S241.INIT=16'h9996;
  LUT4 ZFF_Y1_10_rep1_RNI41DU(.I0(ZFF_Y1_15_rep1),.I1(ZFF_Y1_16_rep1),.I2(un9_11_22_rep1),.I3(un9_11_23_rep1),.O(un9_6_0_axb_16));
defparam ZFF_Y1_10_rep1_RNI41DU.INIT=16'h9C63;
  LUT4 ZFF_Y1_17_rep1_RNINTFL(.I0(ZFF_Y1_16_rep1),.I1(ZFF_Y1_17_rep1),.I2(un9_10[8:8]),.I3(un9_11_23_rep1),.O(un9_6_0_axb_17));
defparam ZFF_Y1_17_rep1_RNINTFL.INIT=16'h96C3;
  LUT3 desc131(.I0(ZFF_Y1[17:17]),.I1(un9_8[6:6]),.I2(un9_10[8:8]),.O(un9_6_0_axb_18));
defparam desc131.INIT=8'hC9;
  LUT4 desc132(.I0(ZFF_Y1[17:17]),.I1(un9_8[6:6]),.I2(un9_8[7:7]),.I3(un9_11_23_rep1),.O(un9_6_0_axb_19));
defparam desc132.INIT=16'h4BB4;
  LUT4 ZFF_Y1_11_rep1_RNI5DD51(.I0(ZFF_Y1[3:3]),.I1(ZFF_Y1_15_rep1),.I2(un9_8[7:7]),.I3(un9_11_23_rep1),.O(un9_6_0_axb_20));
defparam ZFF_Y1_11_rep1_RNI5DD51.INIT=16'h9666;
  LUT4 un9_11_s_10_RNIOI0N1(.I0(ZFF_Y1[15:15]),.I1(un9_11[26:26]),.I2(un9_11[31:31]),.I3(un9_11[32:32]),.O(un9_6_0_axb_32));
defparam un9_11_s_10_RNIOI0N1.INIT=16'h956A;
  LUT4 un9_11_s_11_RNISK0N1(.I0(ZFF_Y1[15:15]),.I1(ZFF_Y1[16:16]),.I2(un9_11[32:32]),.I3(un9_11[33:33]),.O(un9_6_0_axb_33));
defparam un9_11_s_11_RNISK0N1.INIT=16'h936C;
  LUT4 un9_11_s_12_RNI0N0N1(.I0(ZFF_Y1[16:16]),.I1(ZFF_Y1[17:17]),.I2(un9_11[33:33]),.I3(un9_11[34:34]),.O(un9_6_0_axb_34));
defparam un9_11_s_12_RNI0N0N1.INIT=16'h936C;
  LUT3 un9_11_s_13_RNIKNH81(.I0(ZFF_Y1[17:17]),.I1(un9_11[34:34]),.I2(un9_11[35:35]),.O(un9_6_0_axb_35));
defparam un9_11_s_13_RNIKNH81.INIT=8'hD2;
  LUT3 un9_11_s_15_RNIMNH81(.I0(ZFF_Y1[17:17]),.I1(un9_11[35:35]),.I2(un9_11[36:36]),.O(un9_6_0_axb_36));
defparam un9_11_s_15_RNIMNH81.INIT=8'h78;
  LUT2 un9_6_0_axb_37_cZ(.I0(ZFF_Y1[17:17]),.I1(un9_11[37:37]),.O(un9_6_0_axb_37));
defparam un9_6_0_axb_37_cZ.INIT=4'h6;
  LUT1 un9_6_0_axb_38_cZ(.I0(un9_11[38:38]),.O(un9_6_0_axb_38));
defparam un9_6_0_axb_38_cZ.INIT=2'h2;
  LUT1 un9_6_0_axb_39_cZ(.I0(un9_11[39:39]),.O(un9_6_0_axb_39));
defparam un9_6_0_axb_39_cZ.INIT=2'h2;
  LUT2 un9_6_0_axb_40_cZ(.I0(ZFF_Y1[17:17]),.I1(un9_11[40:40]),.O(un9_6_0_axb_40));
defparam un9_6_0_axb_40_cZ.INIT=4'h6;
  LUT2 un9_6_0_axb_41_cZ(.I0(ZFF_Y1[17:17]),.I1(un9_11[41:41]),.O(un9_6_0_axb_41));
defparam un9_6_0_axb_41_cZ.INIT=4'h6;
  LUT1 un9_6_0_axb_42_cZ(.I0(un9_11[42:42]),.O(un9_6_0_axb_42));
defparam un9_6_0_axb_42_cZ.INIT=2'h2;
  LUT2 un9_6_0_axb_43_cZ(.I0(ZFF_Y1[17:17]),.I1(un9_11[43:43]),.O(un9_6_0_axb_43));
defparam un9_6_0_axb_43_cZ.INIT=4'h6;
  LUT1 un9_6_0_axb_44_cZ(.I0(un9_11[44:44]),.O(un9_6_0_axb_44));
defparam un9_6_0_axb_44_cZ.INIT=2'h2;
  LUT2 un9_6_0_axb_45_cZ(.I0(ZFF_Y1[17:17]),.I1(un9_11[45:45]),.O(un9_6_0_axb_45));
defparam un9_6_0_axb_45_cZ.INIT=4'h6;
  LUT1 un9_6_0_axb_46_cZ(.I0(un9_11[46:46]),.O(un9_6_0_axb_46));
defparam un9_6_0_axb_46_cZ.INIT=2'h2;
  LUT2 un9_8_cry_0_RNO_cZ(.I0(ZFF_Y1_3_rep1),.I1(ZFF_Y1_6_rep1),.O(un9_8_cry_0_RNO));
defparam un9_8_cry_0_RNO_cZ.INIT=4'h9;
  LUT2 un9_8_axb_1_cZ(.I0(ZFF_Y1_4_rep1),.I1(un9_8_6_rep1),.O(un9_8_axb_1));
defparam un9_8_axb_1_cZ.INIT=4'h6;
  LUT2 un9_8_axb_2_cZ(.I0(ZFF_Y1_8_rep1),.I1(un9_8_7_rep1),.O(un9_8_axb_2));
defparam un9_8_axb_2_cZ.INIT=4'h9;
  LUT2 un9_8_axb_3_cZ(.I0(ZFF_Y1_3_rep1),.I1(ZFF_Y1_fast[9:9]),.O(un9_8_axb_3));
defparam un9_8_axb_3_cZ.INIT=4'h9;
  LUT2 un9_8_axb_4_cZ(.I0(ZFF_Y1_7_rep1),.I1(un9_11_22_rep1),.O(un9_8_axb_4));
defparam un9_8_axb_4_cZ.INIT=4'h9;
  LUT3 un9_8_axb_5_cZ(.I0(ZFF_Y1_fast[8:8]),.I1(un9_8_fast[6:6]),.I2(un9_11_fast[23:23]),.O(un9_8_axb_5));
defparam un9_8_axb_5_cZ.INIT=8'h69;
  LUT4 desc133(.I0(ZFF_Y1_fast[6:6]),.I1(ZFF_Y1_fast[8:8]),.I2(un9_8_fast[6:6]),.I3(un9_10_8_rep1),.O(un9_8_axb_6));
defparam desc133.INIT=16'h956A;
  LUT4 un9_8_axb_15_cZ(.I0(ZFF_Y1_9_rep1),.I1(ZFF_Y1_fast[8:8]),.I2(un9_8_6_rep1),.I3(un9_8_7_rep1),.O(un9_8_axb_15));
defparam un9_8_axb_15_cZ.INIT=16'hA659;
  LUT4 un9_8_axb_16_cZ(.I0(ZFF_Y1[3:3]),.I1(ZFF_Y1_9_rep1),.I2(un9_8_7_rep1),.I3(un9_11_22_rep1),.O(un9_8_axb_16));
defparam un9_8_axb_16_cZ.INIT=16'hA659;
  LUT4 un9_8_axb_19_cZ(.I0(ZFF_Y1_5_rep1),.I1(ZFF_Y1_6_rep1),.I2(un9_11_25_rep1),.I3(un9_11_fast[24:24]),.O(un9_8_axb_19));
defparam un9_8_axb_19_cZ.INIT=16'h96C3;
  LUT4 un9_8_axb_20_cZ(.I0(ZFF_Y1[7:7]),.I1(ZFF_Y1_6_rep1),.I2(un9_11_25_rep1),.I3(un9_11_26_rep1),.O(un9_8_axb_20));
defparam un9_8_axb_20_cZ.INIT=16'h9A65;
  LUT4 desc134(.I0(ZFF_Y1[7:7]),.I1(ZFF_Y1[8:8]),.I2(ZFF_Y1_15_rep1),.I3(un9_11[26:26]),.O(un9_8_axb_21));
defparam desc134.INIT=16'h693C;
  LUT4 desc135(.I0(ZFF_Y1[8:8]),.I1(ZFF_Y1[9:9]),.I2(ZFF_Y1_15_rep1),.I3(ZFF_Y1_16_rep1),.O(un9_8_axb_22));
defparam desc135.INIT=16'hC639;
  LUT3 desc136(.I0(ZFF_Y1[9:9]),.I1(ZFF_Y1_16_rep1),.I2(un9_11[22:22]),.O(un9_8_axb_23));
defparam desc136.INIT=8'h2D;
  LUT2 un9_8_axb_24_cZ(.I0(un9_11[22:22]),.I1(un9_11[23:23]),.O(un9_8_axb_24));
defparam un9_8_axb_24_cZ.INIT=4'h9;
  LUT2 un9_8_axb_25_cZ(.I0(un9_11[23:23]),.I1(un9_11[24:24]),.O(un9_8_axb_25));
defparam un9_8_axb_25_cZ.INIT=4'h9;
  LUT2 un9_8_axb_26_cZ(.I0(un9_11[24:24]),.I1(un9_11[25:25]),.O(un9_8_axb_26));
defparam un9_8_axb_26_cZ.INIT=4'h9;
  LUT2 un9_8_axb_27_cZ(.I0(un9_11[25:25]),.I1(un9_11[26:26]),.O(un9_8_axb_27));
defparam un9_8_axb_27_cZ.INIT=4'h9;
  LUT2 un9_8_axb_28_cZ(.I0(ZFF_Y1[15:15]),.I1(un9_11[26:26]),.O(un9_8_axb_28));
defparam un9_8_axb_28_cZ.INIT=4'h9;
  LUT1 un9_8_cry_30_RNO_cZ(.I0(ZFF_Y1[16:16]),.O(un9_8_cry_30_RNO));
defparam un9_8_cry_30_RNO_cZ.INIT=2'h1;
  LUT1 un9_10_axb_1_cZ(.I0(ZFF_Y1_3_rep1),.O(un9_10_axb_1));
defparam un9_10_axb_1_cZ.INIT=2'h2;
  LUT3 un9_10_axb_2_cZ(.I0(ZFF_Y1_4_rep1),.I1(ZFF_Y1_fast[9:9]),.I2(un9_8_7_rep1),.O(un9_10_axb_2));
defparam un9_10_axb_2_cZ.INIT=8'h96;
  LUT4 ZFF_Y1_8_rep1_RNIATJ91(.I0(ZFF_Y1_3_rep1),.I1(ZFF_Y1_4_rep1),.I2(ZFF_Y1_7_rep1),.I3(ZFF_Y1_8_rep1),.O(un9_10_axb_4));
defparam ZFF_Y1_8_rep1_RNIATJ91.INIT=16'h936C;
  LUT4 desc137(.I0(ZFF_Y1[15:15]),.I1(un9_11[23:23]),.I2(un9_11[24:24]),.I3(un9_11[26:26]),.O(un9_10_axb_25));
defparam desc137.INIT=16'h965A;
  LUT4 desc138(.I0(ZFF_Y1[15:15]),.I1(ZFF_Y1[16:16]),.I2(un9_11[24:24]),.I3(un9_11[25:25]),.O(un9_10_axb_26));
defparam desc138.INIT=16'h936C;
  LUT3 desc139(.I0(ZFF_Y1[16:16]),.I1(un9_11[25:25]),.I2(un9_11[26:26]),.O(un9_10_axb_27));
defparam desc139.INIT=8'h78;
  LUT1 un9_10_axb_28_cZ(.I0(ZFF_Y1[15:15]),.O(un9_10_axb_28));
defparam un9_10_axb_28_cZ.INIT=2'h2;
  LUT1 un9_10_axb_29_cZ(.I0(ZFF_Y1[16:16]),.O(un9_10_axb_29));
defparam un9_10_axb_29_cZ.INIT=2'h2;
  LUT4 un10_axb_3_cZ(.I0(ZFF_Y2[1:1]),.I1(ZFF_Y2[3:3]),.I2(ZFF_Y2[7:7]),.I3(un10_6[9:9]),.O(un10_axb_3));
defparam un10_axb_3_cZ.INIT=16'h9C63;
  LUT3 un10_axb_6_cZ(.I0(un10_10),.I1(ZFF_Y2[6:6]),.I2(un10_6[12:12]),.O(un10_axb_6));
defparam un10_axb_6_cZ.INIT=8'h69;
  LUT4 un10_axb_7_cZ(.I0(un10_10),.I1(ZFF_Y2[6:6]),.I2(ZFF_Y2[7:7]),.I3(un10_6[13:13]),.O(un10_axb_7));
defparam un10_axb_7_cZ.INIT=16'hD22D;
  LUT3 un10_axb_8_cZ(.I0(ZFF_Y2[6:6]),.I1(ZFF_Y2[14:14]),.I2(un10_6[14:14]),.O(un10_axb_8));
defparam un10_axb_8_cZ.INIT=8'h96;
  LUT4 un10_axb_24_cZ(.I0(un10_6[29:29]),.I1(un10_6[30:30]),.I2(un10_8[29:29]),.I3(un10_8[30:30]),.O(un10_axb_24));
defparam un10_axb_24_cZ.INIT=16'h36C9;
  LUT4 un10_axb_25_cZ(.I0(un10_6[30:30]),.I1(un10_6[31:31]),.I2(un10_8[30:30]),.I3(un10_8[31:31]),.O(un10_axb_25));
defparam un10_axb_25_cZ.INIT=16'h36C9;
  LUT4 un10_axb_26_cZ(.I0(un10_6[31:31]),.I1(un10_6[32:32]),.I2(un10_8[31:31]),.I3(un10_8[32:32]),.O(un10_axb_26));
defparam un10_axb_26_cZ.INIT=16'h36C9;
  LUT4 un10_axb_27_cZ(.I0(un10_6[32:32]),.I1(un10_6[33:33]),.I2(un10_8[32:32]),.I3(un10_8[33:33]),.O(un10_axb_27));
defparam un10_axb_27_cZ.INIT=16'h36C9;
  LUT4 un10_axb_28_cZ(.I0(un10_6[33:33]),.I1(un10_6[34:34]),.I2(un10_8[33:33]),.I3(un10_8[34:34]),.O(un10_axb_28));
defparam un10_axb_28_cZ.INIT=16'h36C9;
  LUT4 un10_6_s_25_RNIAK6M1(.I0(un10_6[34:34]),.I1(un10_6[35:35]),.I2(un10_8[34:34]),.I3(un10_8[35:35]),.O(un10_axb_29));
defparam un10_6_s_25_RNIAK6M1.INIT=16'hC936;
  LUT4 un10_6_cry_26_outext_RNIGU5L1(.I0(un10_6[35:35]),.I1(un10_6[36:36]),.I2(un10_8[35:35]),.I3(un10_8[36:36]),.O(un10_axb_30));
defparam un10_6_cry_26_outext_RNIGU5L1.INIT=16'h6C93;
  LUT3 un10_6_cry_26_outext_RNI0EU91(.I0(un10_6[36:36]),.I1(un10_8[36:36]),.I2(un10_8[37:37]),.O(un10_axb_31));
defparam un10_6_cry_26_outext_RNI0EU91.INIT=8'hE1;
  LUT2 un10_axb_32_cZ(.I0(un10_8[37:37]),.I1(un10_8[38:38]),.O(un10_axb_32));
defparam un10_axb_32_cZ.INIT=4'h9;
  LUT2 un10_axb_33_cZ(.I0(un10_8[38:38]),.I1(un10_8[39:39]),.O(un10_axb_33));
defparam un10_axb_33_cZ.INIT=4'h9;
  LUT2 un10_axb_34_cZ(.I0(un10_8[39:39]),.I1(un10_8[40:40]),.O(un10_axb_34));
defparam un10_axb_34_cZ.INIT=4'h9;
  LUT2 un10_axb_35_cZ(.I0(un10_8[40:40]),.I1(un10_8[41:41]),.O(un10_axb_35));
defparam un10_axb_35_cZ.INIT=4'h9;
  LUT2 un10_axb_36_cZ(.I0(un10_8[41:41]),.I1(un10_8[42:42]),.O(un10_axb_36));
defparam un10_axb_36_cZ.INIT=4'h9;
  LUT2 un10_axb_37_cZ(.I0(un10_8[42:42]),.I1(un10_8[43:43]),.O(un10_axb_37));
defparam un10_axb_37_cZ.INIT=4'h6;
  LUT1 desc140(.I0(un10_8[44:44]),.O(un10_8_i[44:44]));
defparam desc140.INIT=2'h1;
  LUT1 desc141(.I0(un10_8[45:45]),.O(un10_8_i[45:45]));
defparam desc141.INIT=2'h1;
  LUT1 un10_8_s_28_RNIMQRF(.I0(un10_8[47:47]),.O(un10_cry_40_sf));
defparam un10_8_s_28_RNIMQRF.INIT=2'h1;
  LUT4 desc142(.I0(ZFF_Y2[1:1]),.I1(ZFF_Y2[2:2]),.I2(ZFF_Y2[9:9]),.I3(ZFF_Y2[10:10]),.O(un10_6_axb_1));
defparam desc142.INIT=16'h9C63;
  LUT4 desc143(.I0(ZFF_Y2[2:2]),.I1(ZFF_Y2[3:3]),.I2(ZFF_Y2[10:10]),.I3(ZFF_Y2[11:11]),.O(un10_6_axb_2));
defparam desc143.INIT=16'h9C63;
  LUT4 desc144(.I0(ZFF_Y2[11:11]),.I1(ZFF_Y2[12:12]),.I2(ZFF_Y2[15:15]),.I3(ZFF_Y2[16:16]),.O(un10_6_axb_21));
defparam desc144.INIT=16'hC639;
  LUT4 desc145(.I0(ZFF_Y2[12:12]),.I1(ZFF_Y2[13:13]),.I2(ZFF_Y2[16:16]),.I3(ZFF_Y2[17:17]),.O(un10_6_axb_22));
defparam desc145.INIT=16'hC639;
  LUT3 desc146(.I0(ZFF_Y2[13:13]),.I1(ZFF_Y2[14:14]),.I2(ZFF_Y2[17:17]),.O(un10_6_axb_23));
defparam desc146.INIT=8'hC9;
  LUT3 desc147(.I0(ZFF_Y2[14:14]),.I1(ZFF_Y2[15:15]),.I2(ZFF_Y2[17:17]),.O(un10_6_axb_24));
defparam desc147.INIT=8'hC9;
  LUT3 desc148(.I0(ZFF_Y2[15:15]),.I1(ZFF_Y2[16:16]),.I2(ZFF_Y2[17:17]),.O(un10_6_axb_25));
defparam desc148.INIT=8'hC9;
  LUT2 desc149(.I0(ZFF_Y2[16:16]),.I1(ZFF_Y2[17:17]),.O(un10_6_axb_26));
defparam desc149.INIT=4'h2;
  LUT1 un8_0_0_cry_0_RNO(.I0(ZFF_X2[0:0]),.O(N_3207_i));
defparam un8_0_0_cry_0_RNO.INIT=2'h1;
  LUT1 un8_0_0_cry_1_RNO(.I0(ZFF_X2[1:1]),.O(N_3204_i));
defparam un8_0_0_cry_1_RNO.INIT=2'h1;
  LUT1 un8_0_0_cry_2_RNO(.I0(ZFF_X2[2:2]),.O(N_3201_i));
defparam un8_0_0_cry_2_RNO.INIT=2'h1;
  LUT1 un8_0_0_cry_3_RNO(.I0(ZFF_X2[3:3]),.O(N_3198_i));
defparam un8_0_0_cry_3_RNO.INIT=2'h1;
  LUT1 un8_0_0_cry_4_RNO(.I0(ZFF_X2[4:4]),.O(N_3195_i));
defparam un8_0_0_cry_4_RNO.INIT=2'h1;
  LUT2 un8_0_0_cry_5_RNO(.I0(ZFF_X2[0:0]),.I1(ZFF_X2[5:5]),.O(un8_0_6[5:5]));
defparam un8_0_0_cry_5_RNO.INIT=4'h9;
  LUT1 un8_0_0_cry_6_RNO(.I0(un8_0_6[6:6]),.O(un8_0_0_cry_6_sf));
defparam un8_0_0_cry_6_RNO.INIT=2'h2;
  LUT2 un8_0_0_axb_7_cZ(.I0(ZFF_X2[2:2]),.I1(un8_0_6[7:7]),.O(un8_0_0_axb_7));
defparam un8_0_0_axb_7_cZ.INIT=4'h6;
  LUT2 un8_0_0_axb_8_cZ(.I0(ZFF_X2[0:0]),.I1(un8_0_6[8:8]),.O(un8_0_0_axb_8));
defparam un8_0_0_axb_8_cZ.INIT=4'h6;
  LUT2 un8_0_0_axb_9_cZ(.I0(ZFF_X2[1:1]),.I1(un8_0_6[9:9]),.O(un8_0_0_axb_9));
defparam un8_0_0_axb_9_cZ.INIT=4'h6;
  LUT3 un8_0_0_axb_10_cZ(.I0(ZFF_X2[2:2]),.I1(ZFF_X2[3:3]),.I2(un8_0_6[10:10]),.O(un8_0_0_axb_10));
defparam un8_0_0_axb_10_cZ.INIT=8'h96;
  LUT4 un8_0_0_axb_12_cZ(.I0(un8_0_6[11:11]),.I1(un8_0_6[12:12]),.I2(un8_0_8[11:11]),.I3(un8_0_8[12:12]),.O(un8_0_0_axb_12));
defparam un8_0_0_axb_12_cZ.INIT=16'h936C;
  LUT4 un8_0_0_axb_13_cZ(.I0(un8_0_6[12:12]),.I1(un8_0_6[13:13]),.I2(un8_0_8[12:12]),.I3(un8_0_8[13:13]),.O(un8_0_0_axb_13));
defparam un8_0_0_axb_13_cZ.INIT=16'h936C;
  LUT4 un8_0_0_axb_14_cZ(.I0(un8_0_6[13:13]),.I1(un8_0_6[14:14]),.I2(un8_0_8[13:13]),.I3(un8_0_8[14:14]),.O(un8_0_0_axb_14));
defparam un8_0_0_axb_14_cZ.INIT=16'h936C;
  LUT4 un8_0_8_s_20_RNI1AD71(.I0(un8_0_8[29:29]),.I1(un8_0_8[30:30]),.I2(un8_0_9[29:29]),.I3(un8_0_9[30:30]),.O(un8_0_0_axb_30));
defparam un8_0_8_s_20_RNI1AD71.INIT=16'h936C;
  LUT4 un8_0_8_s_20_RNISAD71(.I0(un8_0_8[30:30]),.I1(un8_0_8[31:31]),.I2(un8_0_9[30:30]),.I3(un8_0_9[31:31]),.O(un8_0_0_axb_31));
defparam un8_0_8_s_20_RNISAD71.INIT=16'h936C;
  LUT4 un8_0_8_s_21_RNI0BD71(.I0(un8_0_8[31:31]),.I1(un8_0_8[32:32]),.I2(un8_0_9[31:31]),.I3(un8_0_9[32:32]),.O(un8_0_0_axb_32));
defparam un8_0_8_s_21_RNI0BD71.INIT=16'h936C;
  LUT4 un8_0_8_s_22_RNI4BD71(.I0(un8_0_8[32:32]),.I1(un8_0_8[33:33]),.I2(un8_0_9[32:32]),.I3(un8_0_9[33:33]),.O(un8_0_0_axb_33));
defparam un8_0_8_s_22_RNI4BD71.INIT=16'h936C;
  LUT4 un8_0_8_s_23_RNI8BD71(.I0(un8_0_8[33:33]),.I1(un8_0_8[34:34]),.I2(un8_0_9[33:33]),.I3(un8_0_9[34:34]),.O(un8_0_0_axb_34));
defparam un8_0_8_s_23_RNI8BD71.INIT=16'h936C;
  LUT4 un8_0_8_s_24_RNI3CD71(.I0(un8_0_8[34:34]),.I1(un8_0_8[35:35]),.I2(un8_0_9[34:34]),.I3(un8_0_9[35:35]),.O(un8_0_0_axb_35));
defparam un8_0_8_s_24_RNI3CD71.INIT=16'h936C;
  LUT2 un8_0_6_cry_0_RNO_0(.I0(ZFF_X2[0:0]),.I1(ZFF_X2[5:5]),.O(un8_0_6_cry_0_sf));
defparam un8_0_6_cry_0_RNO_0.INIT=4'h9;
  LUT2 desc150(.I0(ZFF_X2[1:1]),.I1(ZFF_X2[6:6]),.O(un8_0_6_axb_1));
defparam desc150.INIT=4'h9;
  LUT2 desc151(.I0(ZFF_X2[0:0]),.I1(ZFF_X2[7:7]),.O(un8_0_6_axb_2));
defparam desc151.INIT=4'h9;
  LUT3 un8_0_6_axb_3_cZ(.I0(ZFF_X2[1:1]),.I1(ZFF_X2[8:8]),.I2(ZFF_X2_3_rep1),.O(un8_0_6_axb_3));
defparam un8_0_6_axb_3_cZ.INIT=8'h69;
  LUT4 ZFF_X2_14_rep1_RNICVLU(.I0(ZFF_X2[12:12]),.I1(ZFF_X2[13:13]),.I2(ZFF_X2[15:15]),.I3(ZFF_X2_14_rep1),.O(un8_0_6_axb_20));
defparam ZFF_X2_14_rep1_RNICVLU.INIT=16'h963C;
  LUT3 desc152(.I0(ZFF_X2[13:13]),.I1(ZFF_X2[14:14]),.I2(ZFF_X2[15:15]),.O(un8_0_6_axb_21));
defparam desc152.INIT=8'h6C;
  LUT1 un8_0_6_axb_22_cZ(.I0(ZFF_X2[15:15]),.O(un8_0_6_axb_22));
defparam un8_0_6_axb_22_cZ.INIT=2'h2;
  LUT1 un7_0_0_cry_0_thru(.I0(ZFF_X1[0:0]),.O(N_3353_i_0));
defparam un7_0_0_cry_0_thru.INIT=2'h2;
  LUT1 un7_0_0_axb_1_cZ(.I0(ZFF_X1[1:1]),.O(un7_0_0_axb_1));
defparam un7_0_0_axb_1_cZ.INIT=2'h1;
  LUT1 un7_0_0_axb_2_cZ(.I0(ZFF_X1[2:2]),.O(un7_0_0_axb_2));
defparam un7_0_0_axb_2_cZ.INIT=2'h1;
  LUT2 un7_0_0_axb_3_cZ(.I0(ZFF_X1[0:0]),.I1(ZFF_X1[3:3]),.O(un7_0_0_axb_3));
defparam un7_0_0_axb_3_cZ.INIT=4'h9;
  LUT1 un7_0_0_axb_4_cZ(.I0(un7_0_6[4:4]),.O(un7_0_0_axb_4));
defparam un7_0_0_axb_4_cZ.INIT=2'h2;
  LUT1 un7_0_0_axb_5_cZ(.I0(un7_0_6[5:5]),.O(un7_0_0_axb_5));
defparam un7_0_0_axb_5_cZ.INIT=2'h2;
  LUT1 un7_0_0_axb_6_cZ(.I0(un7_0_6[6:6]),.O(un7_0_0_axb_6));
defparam un7_0_0_axb_6_cZ.INIT=2'h2;
  LUT1 un7_0_0_axb_7_cZ(.I0(un7_0_6[7:7]),.O(un7_0_0_axb_7));
defparam un7_0_0_axb_7_cZ.INIT=2'h2;
  LUT2 un7_0_0_axb_8_cZ(.I0(ZFF_X1[5:5]),.I1(un7_0_6[8:8]),.O(un7_0_0_axb_8));
defparam un7_0_0_axb_8_cZ.INIT=4'h6;
  LUT3 un7_0_0_cry_9_RNO(.I0(ZFF_X1[0:0]),.I1(ZFF_X1[3:3]),.I2(un7_0_6[9:9]),.O(un7_0_0_axb_9));
defparam un7_0_0_cry_9_RNO.INIT=8'h96;
  LUT4 un7_0_0_axb_18_cZ(.I0(un7_0_0_o5_17),.I1(un7_0_6[18:18]),.I2(un7_0_8[18:18]),.I3(un7_0_10[18:18]),.O(un7_0_0_axb_18));
defparam un7_0_0_axb_18_cZ.INIT=16'h6996;
  LUT4 un7_0_10_s_17_RNIKBU01(.I0(un7_0_8[34:34]),.I1(un7_0_8[35:35]),.I2(un7_0_10[34:34]),.I3(un7_0_10[35:35]),.O(un7_0_0_axb_35));
defparam un7_0_10_s_17_RNIKBU01.INIT=16'h936C;
  LUT4 un7_0_10_s_17_RNIOBU01(.I0(un7_0_8[35:35]),.I1(un7_0_8[36:36]),.I2(un7_0_10[35:35]),.I3(un7_0_10[36:36]),.O(un7_0_0_axb_36));
defparam un7_0_10_s_17_RNIOBU01.INIT=16'h936C;
  LUT4 un7_0_10_s_18_RNISBU01(.I0(un7_0_8[36:36]),.I1(un7_0_8[37:37]),.I2(un7_0_10[36:36]),.I3(un7_0_10[37:37]),.O(un7_0_0_axb_37));
defparam un7_0_10_s_18_RNISBU01.INIT=16'h936C;
  LUT4 un7_0_10_s_20_RNI4VV9(.I0(ZFF_X1[16:16]),.I1(un7_0_8[38:38]),.I2(un7_0_10[38:38]),.I3(un7_0_10[39:39]),.O(un7_0_0_axb_39));
defparam un7_0_10_s_20_RNI4VV9.INIT=16'hBD42;
  LUT3 un7_0_10_s_22_RNI88V5(.I0(ZFF_X1[16:16]),.I1(un7_0_10[39:39]),.I2(un7_0_10[40:40]),.O(un7_0_0_axb_40));
defparam un7_0_10_s_22_RNI88V5.INIT=8'hD2;
  LUT3 un7_0_10_s_23_RNIA8V5(.I0(ZFF_X1[16:16]),.I1(un7_0_10[40:40]),.I2(un7_0_10[41:41]),.O(un7_0_0_axb_41));
defparam un7_0_10_s_23_RNIA8V5.INIT=8'h78;
  LUT1 un7_0_0_axb_42_cZ(.I0(un7_0_10[42:42]),.O(un7_0_0_axb_42));
defparam un7_0_0_axb_42_cZ.INIT=2'h2;
  LUT1 un7_0_0_axb_43_cZ(.I0(un7_0_10[43:43]),.O(un7_0_0_axb_43));
defparam un7_0_0_axb_43_cZ.INIT=2'h2;
  LUT2 un7_0_0_axb_44_cZ(.I0(ZFF_X1[16:16]),.I1(un7_0_10[44:44]),.O(un7_0_0_axb_44));
defparam un7_0_0_axb_44_cZ.INIT=4'h6;
  LUT2 un7_0_6_cry_0_RNO(.I0(ZFF_X1_0_rep1),.I1(ZFF_X1_3_rep1),.O(un7_0_6[3:3]));
defparam un7_0_6_cry_0_RNO.INIT=4'h9;
  LUT2 desc153(.I0(ZFF_X1_fast[1:1]),.I1(ZFF_X1_fast[4:4]),.O(un7_0_6_axb_1));
defparam desc153.INIT=4'h9;
  LUT2 ZFF_X1_2_rep1_RNIFQO1(.I0(ZFF_X1_2_rep1),.I1(ZFF_X1_5_rep1),.O(un7_0_6_axb_2));
defparam ZFF_X1_2_rep1_RNIFQO1.INIT=4'h9;
  LUT3 un7_0_6_axb_3_cZ(.I0(ZFF_X1_fast[0:0]),.I1(ZFF_X1_fast[3:3]),.I2(ZFF_X1_fast[6:6]),.O(un7_0_6_axb_3));
defparam un7_0_6_axb_3_cZ.INIT=8'h69;
  LUT4 desc154(.I0(ZFF_X1_9_rep1),.I1(ZFF_X1_fast[2:2]),.I2(ZFF_X1_fast[6:6]),.I3(ZFF_X1_fast[8:8]),.O(un7_0_6_axb_6));
defparam desc154.INIT=16'hA569;
  LUT4 desc155(.I0(ZFF_X1_0_rep1),.I1(ZFF_X1_9_rep1),.I2(ZFF_X1_fast[6:6]),.I3(ZFF_X1_fast[10:10]),.O(un7_0_6_axb_7));
defparam desc155.INIT=16'h9A65;
  LUT4 desc156(.I0(ZFF_X1_0_rep1),.I1(ZFF_X1_fast[1:1]),.I2(ZFF_X1_fast[10:10]),.I3(ZFF_X1_fast[11:11]),.O(un7_0_6_axb_8));
defparam desc156.INIT=16'hC639;
  LUT4 un7_0_6_axb_17_cZ(.I0(ZFF_X1_2_rep1),.I1(ZFF_X1_3_rep1),.I2(ZFF_X1_9_rep1),.I3(ZFF_X1_10_rep1),.O(un7_0_6_axb_17));
defparam un7_0_6_axb_17_cZ.INIT=16'hC639;
  LUT4 un7_0_6_axb_18_cZ(.I0(ZFF_X1[4:4]),.I1(ZFF_X1_3_rep1),.I2(ZFF_X1_10_rep1),.I3(ZFF_X1_11_rep1),.O(un7_0_6_axb_18));
defparam un7_0_6_axb_18_cZ.INIT=16'hA659;
  LUT4 un7_0_6_axb_19_cZ(.I0(ZFF_X1[4:4]),.I1(ZFF_X1_5_rep1),.I2(ZFF_X1_11_rep1),.I3(ZFF_X1_12_rep1),.O(un7_0_6_axb_19));
defparam un7_0_6_axb_19_cZ.INIT=16'hC639;
  LUT4 un7_0_6_axb_20_cZ(.I0(ZFF_X1_5_rep1),.I1(ZFF_X1_6_rep1),.I2(ZFF_X1_12_rep1),.I3(ZFF_X1_13_rep1),.O(un7_0_6_axb_20));
defparam un7_0_6_axb_20_cZ.INIT=16'hC639;
  LUT4 un7_0_6_axb_21_cZ(.I0(ZFF_X1[6:6]),.I1(ZFF_X1[14:14]),.I2(ZFF_X1_7_rep1),.I3(ZFF_X1_13_rep1),.O(un7_0_6_axb_21));
defparam un7_0_6_axb_21_cZ.INIT=16'hC369;
  LUT4 ZFF_X1_7_rep1_RNIC4IV(.I0(ZFF_X1[14:14]),.I1(ZFF_X1_7_rep1),.I2(ZFF_X1_8_rep1),.I3(ZFF_X1_15_rep1),.O(un7_0_6_axb_22));
defparam ZFF_X1_7_rep1_RNIC4IV.INIT=16'h4BB4;
  LUT3 ZFF_X1_15_rep1_RNI5UAT(.I0(ZFF_X1[9:9]),.I1(ZFF_X1_8_rep1),.I2(ZFF_X1_15_rep1),.O(un7_0_6_axb_23));
defparam ZFF_X1_15_rep1_RNI5UAT.INIT=8'h65;
  LUT2 desc157(.I0(ZFF_X1[10:10]),.I1(ZFF_X1[16:16]),.O(un7_0_6_axb_24));
defparam desc157.INIT=4'h9;
  LUT1 un7_0_6_axb_25_cZ(.I0(ZFF_X1[11:11]),.O(un7_0_6_axb_25));
defparam un7_0_6_axb_25_cZ.INIT=2'h1;
  LUT1 un7_0_6_axb_26_cZ(.I0(ZFF_X1[12:12]),.O(un7_0_6_axb_26));
defparam un7_0_6_axb_26_cZ.INIT=2'h1;
  LUT1 un7_0_6_axb_27_cZ(.I0(ZFF_X1[13:13]),.O(un7_0_6_axb_27));
defparam un7_0_6_axb_27_cZ.INIT=2'h1;
  LUT1 un7_0_6_axb_28_cZ(.I0(ZFF_X1[14:14]),.O(un7_0_6_axb_28));
defparam un7_0_6_axb_28_cZ.INIT=2'h1;
  LUT1 un7_0_6_axb_29_cZ(.I0(ZFF_X1[15:15]),.O(un7_0_6_axb_29));
defparam un7_0_6_axb_29_cZ.INIT=2'h1;
  LUT2 un7_0_8_axb_1_cZ(.I0(ZFF_X1_4_rep1),.I1(ZFF_X1_7_rep1),.O(un7_0_8_axb_1));
defparam un7_0_8_axb_1_cZ.INIT=4'h6;
  LUT2 un7_0_8_axb_2_cZ(.I0(ZFF_X1_5_rep1),.I1(ZFF_X1_8_rep1),.O(un7_0_8_axb_2));
defparam un7_0_8_axb_2_cZ.INIT=4'h6;
  LUT2 un7_0_8_axb_3_cZ(.I0(ZFF_X1[0:0]),.I1(ZFF_X1_9_rep1),.O(un7_0_8_axb_3));
defparam un7_0_8_axb_3_cZ.INIT=4'h6;
  LUT2 un7_0_8_axb_4_cZ(.I0(ZFF_X1[1:1]),.I1(ZFF_X1_10_rep1),.O(un7_0_8_axb_4));
defparam un7_0_8_axb_4_cZ.INIT=4'h6;
  LUT3 un7_0_8_axb_5_cZ(.I0(ZFF_X1_0_rep1),.I1(ZFF_X1_fast[2:2]),.I2(ZFF_X1_fast[5:5]),.O(un7_0_8_axb_5));
defparam un7_0_8_axb_5_cZ.INIT=8'h96;
  LUT4 ZFF_X1_6_rep1_RNIPNP31(.I0(ZFF_X1[7:7]),.I1(ZFF_X1_6_rep1),.I2(ZFF_X1_15_rep1),.I3(ZFF_X1_fast[14:14]),.O(un7_0_8_axb_20));
defparam ZFF_X1_6_rep1_RNIPNP31.INIT=16'h965A;
  LUT3 desc158(.I0(ZFF_X1[7:7]),.I1(ZFF_X1[8:8]),.I2(ZFF_X1[15:15]),.O(un7_0_8_axb_21));
defparam desc158.INIT=8'h6C;
  LUT1 un7_0_8_axb_22_cZ(.I0(ZFF_X1[9:9]),.O(un7_0_8_axb_22));
defparam un7_0_8_axb_22_cZ.INIT=2'h2;
  LUT1 un7_0_8_axb_23_cZ(.I0(ZFF_X1[10:10]),.O(un7_0_8_axb_23));
defparam un7_0_8_axb_23_cZ.INIT=2'h2;
  LUT1 un7_0_8_axb_24_cZ(.I0(ZFF_X1[11:11]),.O(un7_0_8_axb_24));
defparam un7_0_8_axb_24_cZ.INIT=2'h2;
  LUT1 un7_0_8_axb_25_cZ(.I0(ZFF_X1[12:12]),.O(un7_0_8_axb_25));
defparam un7_0_8_axb_25_cZ.INIT=2'h2;
  LUT1 un7_0_8_axb_26_cZ(.I0(ZFF_X1[13:13]),.O(un7_0_8_axb_26));
defparam un7_0_8_axb_26_cZ.INIT=2'h2;
  LUT1 un7_0_8_axb_27_cZ(.I0(ZFF_X1[14:14]),.O(un7_0_8_axb_27));
defparam un7_0_8_axb_27_cZ.INIT=2'h2;
  LUT1 un7_0_8_axb_28_cZ(.I0(ZFF_X1[15:15]),.O(un7_0_8_axb_28));
defparam un7_0_8_axb_28_cZ.INIT=2'h2;
  LUT2 un6_0_8_axb_0(.I0(ZFF_X0_3_rep1),.I1(ZFF_X0_fast[2:2]),.O(un6_0_8[10:10]));
defparam un6_0_8_axb_0.INIT=4'h6;
  LUT2 un6_0_8_axb_1_cZ(.I0(ZFF_X0_3_rep1),.I1(ZFF_X0_fast[4:4]),.O(un6_0_8_axb_1));
defparam un6_0_8_axb_1_cZ.INIT=4'h6;
  LUT3 un6_0_8_axb_2_cZ(.I0(ZFF_X0_fast[4:4]),.I1(ZFF_X0_fast[5:5]),.I2(ZFF_X0_fast[7:7]),.O(un6_0_8_axb_2));
defparam un6_0_8_axb_2_cZ.INIT=8'h96;
  LUT4 un6_0_8_axb_12_cZ(.I0(ZFF_X0_1_rep1),.I1(ZFF_X0_2_rep1),.I2(ZFF_X0_7_rep1),.I3(ZFF_X0_fast[6:6]),.O(un6_0_8_axb_12));
defparam un6_0_8_axb_12_cZ.INIT=16'h96C3;
  LUT4 un6_0_8_axb_21_cZ(.I0(ZFF_X0[10:10]),.I1(ZFF_X0[11:11]),.I2(ZFF_X0_15_rep1),.I3(ZFF_X0_16_rep1),.O(un6_0_8_axb_21));
defparam un6_0_8_axb_21_cZ.INIT=16'h9C39;
  LUT2 un6_0_8_axb_22_cZ(.I0(ZFF_X0[11:11]),.I1(ZFF_X0[12:12]),.O(un6_0_8_axb_22));
defparam un6_0_8_axb_22_cZ.INIT=4'h9;
  LUT2 un6_0_8_axb_23_cZ(.I0(ZFF_X0[12:12]),.I1(ZFF_X0[13:13]),.O(un6_0_8_axb_23));
defparam un6_0_8_axb_23_cZ.INIT=4'h9;
  LUT2 un6_0_8_axb_24_cZ(.I0(ZFF_X0[13:13]),.I1(ZFF_X0[14:14]),.O(un6_0_8_axb_24));
defparam un6_0_8_axb_24_cZ.INIT=4'h9;
  LUT2 un6_0_8_axb_25_cZ(.I0(ZFF_X0[14:14]),.I1(ZFF_X0[15:15]),.O(un6_0_8_axb_25));
defparam un6_0_8_axb_25_cZ.INIT=4'h9;
  LUT2 un6_0_8_axb_26_cZ(.I0(ZFF_X0[15:15]),.I1(ZFF_X0[16:16]),.O(un6_0_8_axb_26));
defparam un6_0_8_axb_26_cZ.INIT=4'h6;
  LUT2 un8_0_8_axb_0(.I0(ZFF_X2_3_rep1),.I1(ZFF_X2_fast[2:2]),.O(un8_0_8[10:10]));
defparam un8_0_8_axb_0.INIT=4'h6;
  LUT2 un8_0_8_axb_1_cZ(.I0(ZFF_X2_3_rep1),.I1(ZFF_X2_fast[4:4]),.O(un8_0_8_axb_1));
defparam un8_0_8_axb_1_cZ.INIT=4'h6;
  LUT3 un8_0_8_axb_2_cZ(.I0(ZFF_X2_fast[4:4]),.I1(ZFF_X2_fast[5:5]),.I2(ZFF_X2_fast[7:7]),.O(un8_0_8_axb_2));
defparam un8_0_8_axb_2_cZ.INIT=8'h96;
  LUT4 un8_0_8_axb_12_cZ(.I0(ZFF_X2[7:7]),.I1(ZFF_X2_2_rep1),.I2(ZFF_X2_6_rep1),.I3(ZFF_X2_fast[1:1]),.O(un8_0_8_axb_12));
defparam un8_0_8_axb_12_cZ.INIT=16'h9969;
  LUT4 un8_0_8_axb_21_cZ(.I0(ZFF_X2[10:10]),.I1(ZFF_X2[11:11]),.I2(ZFF_X2[16:16]),.I3(ZFF_X2_15_rep1),.O(un8_0_8_axb_21));
defparam un8_0_8_axb_21_cZ.INIT=16'h93C9;
  LUT2 un8_0_8_axb_22_cZ(.I0(ZFF_X2[11:11]),.I1(ZFF_X2[12:12]),.O(un8_0_8_axb_22));
defparam un8_0_8_axb_22_cZ.INIT=4'h9;
  LUT2 un8_0_8_axb_23_cZ(.I0(ZFF_X2[12:12]),.I1(ZFF_X2[13:13]),.O(un8_0_8_axb_23));
defparam un8_0_8_axb_23_cZ.INIT=4'h9;
  LUT2 un8_0_8_axb_24_cZ(.I0(ZFF_X2[13:13]),.I1(ZFF_X2[14:14]),.O(un8_0_8_axb_24));
defparam un8_0_8_axb_24_cZ.INIT=4'h9;
  LUT2 un8_0_8_axb_25_cZ(.I0(ZFF_X2[14:14]),.I1(ZFF_X2[15:15]),.O(un8_0_8_axb_25));
defparam un8_0_8_axb_25_cZ.INIT=4'h9;
  LUT2 un8_0_8_axb_26_cZ(.I0(ZFF_X2[15:15]),.I1(ZFF_X2[16:16]),.O(un8_0_8_axb_26));
defparam un8_0_8_axb_26_cZ.INIT=4'h6;
  LUT2 un10_8_axb_0_cZ(.I0(ZFF_Y2[10:10]),.I1(ZFF_Y2_fast[17:17]),.O(un10_8_axb_0));
defparam un10_8_axb_0_cZ.INIT=4'h9;
  LUT2 un10_8_axb_1_cZ(.I0(ZFF_Y2[11:11]),.I1(ZFF_Y2_fast[17:17]),.O(un10_8_axb_1));
defparam un10_8_axb_1_cZ.INIT=4'h9;
  LUT2 un10_8_axb_2_cZ(.I0(ZFF_Y2[12:12]),.I1(ZFF_Y2_fast[17:17]),.O(un10_8_axb_2));
defparam un10_8_axb_2_cZ.INIT=4'h9;
  LUT2 un10_8_axb_3_cZ(.I0(ZFF_Y2[13:13]),.I1(ZFF_Y2_fast[17:17]),.O(un10_8_axb_3));
defparam un10_8_axb_3_cZ.INIT=4'h9;
  LUT2 un10_8_axb_4_cZ(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2_fast[17:17]),.O(un10_8_axb_4));
defparam un10_8_axb_4_cZ.INIT=4'h9;
  LUT1 un10_8_axb_5_cZ(.I0(ZFF_Y2[0:0]),.O(un10_8_axb_5));
defparam un10_8_axb_5_cZ.INIT=2'h1;
  LUT1 un10_8_axb_6_cZ(.I0(ZFF_Y2[1:1]),.O(un10_8_axb_6));
defparam un10_8_axb_6_cZ.INIT=2'h1;
  LUT1 un10_8_axb_7_cZ(.I0(ZFF_Y2[2:2]),.O(un10_8_axb_7));
defparam un10_8_axb_7_cZ.INIT=2'h1;
  LUT2 un10_8_axb_8_cZ(.I0(ZFF_Y2[0:0]),.I1(ZFF_Y2[3:3]),.O(un10_8_axb_8));
defparam un10_8_axb_8_cZ.INIT=4'h9;
  LUT2 un10_8_axb_9_cZ(.I0(ZFF_Y2[1:1]),.I1(ZFF_Y2[4:4]),.O(un10_8_axb_9));
defparam un10_8_axb_9_cZ.INIT=4'h9;
  LUT3 un10_8_axb_10_cZ(.I0(ZFF_Y2[0:0]),.I1(ZFF_Y2[2:2]),.I2(ZFF_Y2[5:5]),.O(un10_8_axb_10));
defparam un10_8_axb_10_cZ.INIT=8'h69;
  LUT4 un10_8_axb_25_cZ(.I0(ZFF_Y2[14:14]),.I1(ZFF_Y2[15:15]),.I2(ZFF_Y2[16:16]),.I3(ZFF_Y2[17:17]),.O(un10_8_axb_25));
defparam un10_8_axb_25_cZ.INIT=16'h6C36;
  LUT1 un10_8_axb_26_cZ(.I0(ZFF_Y2[16:16]),.O(un10_8_axb_26));
defparam un10_8_axb_26_cZ.INIT=2'h2;
  LUT1 un10_8_axb_27_cZ(.I0(ZFF_Y2[17:17]),.O(un10_8_axb_27));
defparam un10_8_axb_27_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_cry_1_RNO(.I0(pgZFF_X0[1:1]),.O(pgZFF_X0_i[1:1]));
defparam Y_out_double_2_7_cry_1_RNO.INIT=2'h1;
  LUT1 Y_out_double_2_7_axb_2_cZ(.I0(pgZFF_X0[2:2]),.O(Y_out_double_2_7_axb_2));
defparam Y_out_double_2_7_axb_2_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_3_cZ(.I0(pgZFF_X0[3:3]),.O(Y_out_double_2_7_axb_3));
defparam Y_out_double_2_7_axb_3_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_4_cZ(.I0(pgZFF_X0[4:4]),.O(Y_out_double_2_7_axb_4));
defparam Y_out_double_2_7_axb_4_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_5_cZ(.I0(pgZFF_X0[5:5]),.O(Y_out_double_2_7_axb_5));
defparam Y_out_double_2_7_axb_5_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_6_cZ(.I0(pgZFF_X0[6:6]),.O(Y_out_double_2_7_axb_6));
defparam Y_out_double_2_7_axb_6_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_7_cZ(.I0(pgZFF_X0[7:7]),.O(Y_out_double_2_7_axb_7));
defparam Y_out_double_2_7_axb_7_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_8_cZ(.I0(pgZFF_X0[8:8]),.O(Y_out_double_2_7_axb_8));
defparam Y_out_double_2_7_axb_8_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_9_cZ(.I0(pgZFF_X0[9:9]),.O(Y_out_double_2_7_axb_9));
defparam Y_out_double_2_7_axb_9_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_10_cZ(.I0(pgZFF_X0[10:10]),.O(Y_out_double_2_7_axb_10));
defparam Y_out_double_2_7_axb_10_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_11_cZ(.I0(pgZFF_X0[11:11]),.O(Y_out_double_2_7_axb_11));
defparam Y_out_double_2_7_axb_11_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_12_cZ(.I0(pgZFF_X0[12:12]),.O(Y_out_double_2_7_axb_12));
defparam Y_out_double_2_7_axb_12_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_13_cZ(.I0(pgZFF_X0[13:13]),.O(Y_out_double_2_7_axb_13));
defparam Y_out_double_2_7_axb_13_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_14_cZ(.I0(pgZFF_X0[14:14]),.O(Y_out_double_2_7_axb_14));
defparam Y_out_double_2_7_axb_14_cZ.INIT=2'h2;
  LUT1 Y_out_double_2_7_axb_15_cZ(.I0(pgZFF_X0[16:16]),.O(Y_out_double_2_7_axb_15));
defparam Y_out_double_2_7_axb_15_cZ.INIT=2'h2;
  LUT1 un6_0_9_axb_1_cZ(.I0(ZFF_X0[8:8]),.O(un6_0_9_axb_1));
defparam un6_0_9_axb_1_cZ.INIT=2'h2;
  LUT1 un6_0_9_axb_2_cZ(.I0(ZFF_X0[9:9]),.O(un6_0_9_axb_2));
defparam un6_0_9_axb_2_cZ.INIT=2'h2;
  LUT1 un6_0_9_axb_3_cZ(.I0(ZFF_X0_10_rep1),.O(un6_0_9_axb_3));
defparam un6_0_9_axb_3_cZ.INIT=2'h2;
  LUT1 un6_0_9_axb_4_cZ(.I0(ZFF_X0[11:11]),.O(un6_0_9_axb_4));
defparam un6_0_9_axb_4_cZ.INIT=2'h2;
  LUT2 un6_0_9_axb_5_cZ(.I0(ZFF_X0[13:13]),.I1(ZFF_X0_12_rep1),.O(un6_0_9_axb_5));
defparam un6_0_9_axb_5_cZ.INIT=4'h6;
  LUT1 un6_0_9_axb_6_cZ(.I0(ZFF_X0[13:13]),.O(un6_0_9_axb_6));
defparam un6_0_9_axb_6_cZ.INIT=2'h2;
  LUT1 un6_0_9_axb_7_cZ(.I0(ZFF_X0[14:14]),.O(un6_0_9_axb_7));
defparam un6_0_9_axb_7_cZ.INIT=2'h2;
  LUT1 un6_0_9_axb_8_cZ(.I0(ZFF_X0[0:0]),.O(un6_0_9_axb_8));
defparam un6_0_9_axb_8_cZ.INIT=2'h1;
  LUT1 un6_0_9_axb_9_cZ(.I0(ZFF_X0[1:1]),.O(un6_0_9_axb_9));
defparam un6_0_9_axb_9_cZ.INIT=2'h1;
  LUT1 un6_0_9_axb_10_cZ(.I0(ZFF_X0[2:2]),.O(un6_0_9_axb_10));
defparam un6_0_9_axb_10_cZ.INIT=2'h1;
  LUT2 un6_0_9_axb_11_cZ(.I0(ZFF_X0[0:0]),.I1(ZFF_X0[3:3]),.O(un6_0_9_axb_11));
defparam un6_0_9_axb_11_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_12_cZ(.I0(ZFF_X0[1:1]),.I1(ZFF_X0[4:4]),.O(un6_0_9_axb_12));
defparam un6_0_9_axb_12_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_13_cZ(.I0(ZFF_X0[2:2]),.I1(ZFF_X0[5:5]),.O(un6_0_9_axb_13));
defparam un6_0_9_axb_13_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_14_cZ(.I0(ZFF_X0[3:3]),.I1(ZFF_X0[6:6]),.O(un6_0_9_axb_14));
defparam un6_0_9_axb_14_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_15_cZ(.I0(ZFF_X0[4:4]),.I1(ZFF_X0[7:7]),.O(un6_0_9_axb_15));
defparam un6_0_9_axb_15_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_16_cZ(.I0(ZFF_X0[5:5]),.I1(ZFF_X0[8:8]),.O(un6_0_9_axb_16));
defparam un6_0_9_axb_16_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_17_cZ(.I0(ZFF_X0[6:6]),.I1(ZFF_X0[9:9]),.O(un6_0_9_axb_17));
defparam un6_0_9_axb_17_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_18_cZ(.I0(ZFF_X0[7:7]),.I1(ZFF_X0[10:10]),.O(un6_0_9_axb_18));
defparam un6_0_9_axb_18_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_19_cZ(.I0(ZFF_X0[8:8]),.I1(ZFF_X0[11:11]),.O(un6_0_9_axb_19));
defparam un6_0_9_axb_19_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_20_cZ(.I0(ZFF_X0[9:9]),.I1(ZFF_X0[12:12]),.O(un6_0_9_axb_20));
defparam un6_0_9_axb_20_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_21_cZ(.I0(ZFF_X0[10:10]),.I1(ZFF_X0[13:13]),.O(un6_0_9_axb_21));
defparam un6_0_9_axb_21_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_22_cZ(.I0(ZFF_X0[11:11]),.I1(ZFF_X0[14:14]),.O(un6_0_9_axb_22));
defparam un6_0_9_axb_22_cZ.INIT=4'h9;
  LUT2 un6_0_9_axb_23_cZ(.I0(ZFF_X0[12:12]),.I1(ZFF_X0[15:15]),.O(un6_0_9_axb_23));
defparam un6_0_9_axb_23_cZ.INIT=4'h9;
  LUT1 un6_0_9_axb_24_cZ(.I0(ZFF_X0[13:13]),.O(un6_0_9_axb_24));
defparam un6_0_9_axb_24_cZ.INIT=2'h2;
  LUT1 un6_0_9_axb_25_cZ(.I0(ZFF_X0[14:14]),.O(un6_0_9_axb_25));
defparam un6_0_9_axb_25_cZ.INIT=2'h2;
  LUT1 un6_0_9_axb_26_cZ(.I0(ZFF_X0[15:15]),.O(un6_0_9_axb_26));
defparam un6_0_9_axb_26_cZ.INIT=2'h2;
  LUT1 un8_0_9_axb_1_cZ(.I0(ZFF_X2[8:8]),.O(un8_0_9_axb_1));
defparam un8_0_9_axb_1_cZ.INIT=2'h2;
  LUT1 un8_0_9_axb_2_cZ(.I0(ZFF_X2[9:9]),.O(un8_0_9_axb_2));
defparam un8_0_9_axb_2_cZ.INIT=2'h2;
  LUT1 un8_0_9_axb_3_cZ(.I0(ZFF_X2_10_rep1),.O(un8_0_9_axb_3));
defparam un8_0_9_axb_3_cZ.INIT=2'h2;
  LUT1 un8_0_9_axb_4_cZ(.I0(ZFF_X2[11:11]),.O(un8_0_9_axb_4));
defparam un8_0_9_axb_4_cZ.INIT=2'h2;
  LUT2 un8_0_9_axb_5_cZ(.I0(ZFF_X2[12:12]),.I1(ZFF_X2[13:13]),.O(un8_0_9_axb_5));
defparam un8_0_9_axb_5_cZ.INIT=4'h6;
  LUT1 un8_0_9_axb_6_cZ(.I0(ZFF_X2[13:13]),.O(un8_0_9_axb_6));
defparam un8_0_9_axb_6_cZ.INIT=2'h2;
  LUT1 un8_0_9_axb_7_cZ(.I0(ZFF_X2[14:14]),.O(un8_0_9_axb_7));
defparam un8_0_9_axb_7_cZ.INIT=2'h2;
  LUT1 un8_0_9_axb_8_cZ(.I0(ZFF_X2[0:0]),.O(un8_0_9_axb_8));
defparam un8_0_9_axb_8_cZ.INIT=2'h1;
  LUT1 un8_0_9_axb_9_cZ(.I0(ZFF_X2[1:1]),.O(un8_0_9_axb_9));
defparam un8_0_9_axb_9_cZ.INIT=2'h1;
  LUT1 un8_0_9_axb_10_cZ(.I0(ZFF_X2[2:2]),.O(un8_0_9_axb_10));
defparam un8_0_9_axb_10_cZ.INIT=2'h1;
  LUT2 un8_0_9_axb_11_cZ(.I0(ZFF_X2[0:0]),.I1(ZFF_X2[3:3]),.O(un8_0_9_axb_11));
defparam un8_0_9_axb_11_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_12_cZ(.I0(ZFF_X2[1:1]),.I1(ZFF_X2[4:4]),.O(un8_0_9_axb_12));
defparam un8_0_9_axb_12_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_13_cZ(.I0(ZFF_X2[2:2]),.I1(ZFF_X2[5:5]),.O(un8_0_9_axb_13));
defparam un8_0_9_axb_13_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_14_cZ(.I0(ZFF_X2[3:3]),.I1(ZFF_X2[6:6]),.O(un8_0_9_axb_14));
defparam un8_0_9_axb_14_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_15_cZ(.I0(ZFF_X2[4:4]),.I1(ZFF_X2[7:7]),.O(un8_0_9_axb_15));
defparam un8_0_9_axb_15_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_16_cZ(.I0(ZFF_X2[5:5]),.I1(ZFF_X2[8:8]),.O(un8_0_9_axb_16));
defparam un8_0_9_axb_16_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_17_cZ(.I0(ZFF_X2[6:6]),.I1(ZFF_X2[9:9]),.O(un8_0_9_axb_17));
defparam un8_0_9_axb_17_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_18_cZ(.I0(ZFF_X2[7:7]),.I1(ZFF_X2[10:10]),.O(un8_0_9_axb_18));
defparam un8_0_9_axb_18_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_19_cZ(.I0(ZFF_X2[8:8]),.I1(ZFF_X2[11:11]),.O(un8_0_9_axb_19));
defparam un8_0_9_axb_19_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_20_cZ(.I0(ZFF_X2[9:9]),.I1(ZFF_X2[12:12]),.O(un8_0_9_axb_20));
defparam un8_0_9_axb_20_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_21_cZ(.I0(ZFF_X2[10:10]),.I1(ZFF_X2[13:13]),.O(un8_0_9_axb_21));
defparam un8_0_9_axb_21_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_22_cZ(.I0(ZFF_X2[11:11]),.I1(ZFF_X2[14:14]),.O(un8_0_9_axb_22));
defparam un8_0_9_axb_22_cZ.INIT=4'h9;
  LUT2 un8_0_9_axb_23_cZ(.I0(ZFF_X2[12:12]),.I1(ZFF_X2[15:15]),.O(un8_0_9_axb_23));
defparam un8_0_9_axb_23_cZ.INIT=4'h9;
  LUT1 un8_0_9_axb_24_cZ(.I0(ZFF_X2[13:13]),.O(un8_0_9_axb_24));
defparam un8_0_9_axb_24_cZ.INIT=2'h2;
  LUT1 un8_0_9_axb_25_cZ(.I0(ZFF_X2[14:14]),.O(un8_0_9_axb_25));
defparam un8_0_9_axb_25_cZ.INIT=2'h2;
  LUT1 un8_0_9_axb_26_cZ(.I0(ZFF_X2[15:15]),.O(un8_0_9_axb_26));
defparam un8_0_9_axb_26_cZ.INIT=2'h2;
  LUT2 un9_11_cry_6_RNO_cZ(.I0(ZFF_Y1_fast[15:15]),.I1(un9_10_fast[8:8]),.O(un9_11_cry_6_RNO));
defparam un9_11_cry_6_RNO_cZ.INIT=4'h6;
  LUT2 un9_11_axb_7_cZ(.I0(ZFF_Y1_fast[16:16]),.I1(un9_8_fast[6:6]),.O(un9_11_axb_7));
defparam un9_11_axb_7_cZ.INIT=4'h6;
  LUT2 desc159(.I0(un9_8_fast[7:7]),.I1(un9_10_fast[8:8]),.O(un9_11_axb_8));
defparam desc159.INIT=4'h9;
  LUT2 un9_11_axb_9_cZ(.I0(ZFF_Y1_fast[3:3]),.I1(un9_8_fast[6:6]),.O(un9_11_axb_9));
defparam un9_11_axb_9_cZ.INIT=4'h9;
  LUT2 un9_11_axb_10_cZ(.I0(ZFF_Y1_fast[4:4]),.I1(un9_8_fast[7:7]),.O(un9_11_axb_10));
defparam un9_11_axb_10_cZ.INIT=4'h9;
  LUT2 un9_11_axb_11_cZ(.I0(ZFF_Y1_fast[3:3]),.I1(ZFF_Y1_fast[5:5]),.O(un9_11_axb_11));
defparam un9_11_axb_11_cZ.INIT=4'h9;
  LUT2 un9_11_axb_12_cZ(.I0(ZFF_Y1_fast[4:4]),.I1(ZFF_Y1_fast[6:6]),.O(un9_11_axb_12));
defparam un9_11_axb_12_cZ.INIT=4'h9;
  LUT2 un9_11_axb_13_cZ(.I0(ZFF_Y1_fast[5:5]),.I1(ZFF_Y1_fast[7:7]),.O(un9_11_axb_13));
defparam un9_11_axb_13_cZ.INIT=4'h9;
  LUT2 un9_11_axb_14_cZ(.I0(ZFF_Y1_fast[6:6]),.I1(ZFF_Y1_fast[8:8]),.O(un9_11_axb_14));
defparam un9_11_axb_14_cZ.INIT=4'h9;
  LUT2 un9_11_axb_15_cZ(.I0(ZFF_Y1_fast[7:7]),.I1(ZFF_Y1_fast[9:9]),.O(un9_11_axb_15));
defparam un9_11_axb_15_cZ.INIT=4'h9;
  LUT2 desc160(.I0(ZFF_Y1_fast[8:8]),.I1(un9_11_fast[22:22]),.O(un9_11_axb_16));
defparam desc160.INIT=4'h9;
  LUT2 desc161(.I0(ZFF_Y1_fast[9:9]),.I1(un9_11_fast[23:23]),.O(un9_11_axb_17));
defparam desc161.INIT=4'h9;
  LUT2 un9_11_axb_18_cZ(.I0(un9_11_fast[22:22]),.I1(un9_11_fast[24:24]),.O(un9_11_axb_18));
defparam un9_11_axb_18_cZ.INIT=4'h9;
  LUT2 un9_11_axb_19_cZ(.I0(un9_11_23_rep1),.I1(un9_11_25_rep1),.O(un9_11_axb_19));
defparam un9_11_axb_19_cZ.INIT=4'h9;
  LUT2 un9_11_axb_20_cZ(.I0(un9_11_24_rep1),.I1(un9_11_26_rep1),.O(un9_11_axb_20));
defparam un9_11_axb_20_cZ.INIT=4'h9;
  LUT2 un9_11_axb_21_cZ(.I0(ZFF_Y1_15_rep1),.I1(un9_11_25_rep1),.O(un9_11_axb_21));
defparam un9_11_axb_21_cZ.INIT=4'h9;
  LUT2 un9_11_axb_22_cZ(.I0(ZFF_Y1_16_rep1),.I1(un9_11_26_rep1),.O(un9_11_axb_22));
defparam un9_11_axb_22_cZ.INIT=4'h9;
  LUT1 un9_11_axb_23_cZ(.I0(ZFF_Y1[15:15]),.O(un9_11_axb_23));
defparam un9_11_axb_23_cZ.INIT=2'h1;
  LUT1 un9_11_axb_24_cZ(.I0(ZFF_Y1[16:16]),.O(un9_11_axb_24));
defparam un9_11_axb_24_cZ.INIT=2'h1;
  LUT2 Y_out_double_2_4_axb_1_cZ(.I0(pgZFF_X0[1:1]),.I1(pgZFF_X2[1:1]),.O(Y_out_double_2_4_axb_1));
defparam Y_out_double_2_4_axb_1_cZ.INIT=4'h9;
  LUT2 Y_out_double_2_4_axb_2_cZ(.I0(Y_out_double_2_7[2:2]),.I1(pgZFF_X2[2:2]),.O(Y_out_double_2_4_axb_2));
defparam Y_out_double_2_4_axb_2_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_3_cZ(.I0(Y_out_double_2_7[3:3]),.I1(pgZFF_X2[3:3]),.O(Y_out_double_2_4_axb_3));
defparam Y_out_double_2_4_axb_3_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_4_cZ(.I0(Y_out_double_2_7[4:4]),.I1(pgZFF_X2[4:4]),.O(Y_out_double_2_4_axb_4));
defparam Y_out_double_2_4_axb_4_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_5_cZ(.I0(Y_out_double_2_7[5:5]),.I1(pgZFF_X2[5:5]),.O(Y_out_double_2_4_axb_5));
defparam Y_out_double_2_4_axb_5_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_6_cZ(.I0(Y_out_double_2_7[6:6]),.I1(pgZFF_X2[6:6]),.O(Y_out_double_2_4_axb_6));
defparam Y_out_double_2_4_axb_6_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_7_cZ(.I0(Y_out_double_2_7[7:7]),.I1(pgZFF_X2[7:7]),.O(Y_out_double_2_4_axb_7));
defparam Y_out_double_2_4_axb_7_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_8_cZ(.I0(Y_out_double_2_7[8:8]),.I1(pgZFF_X2[8:8]),.O(Y_out_double_2_4_axb_8));
defparam Y_out_double_2_4_axb_8_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_9_cZ(.I0(Y_out_double_2_7[9:9]),.I1(pgZFF_X2[9:9]),.O(Y_out_double_2_4_axb_9));
defparam Y_out_double_2_4_axb_9_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_10_cZ(.I0(Y_out_double_2_7[10:10]),.I1(pgZFF_X2[10:10]),.O(Y_out_double_2_4_axb_10));
defparam Y_out_double_2_4_axb_10_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_11_cZ(.I0(Y_out_double_2_7[11:11]),.I1(pgZFF_X2[11:11]),.O(Y_out_double_2_4_axb_11));
defparam Y_out_double_2_4_axb_11_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_12_cZ(.I0(Y_out_double_2_7[12:12]),.I1(pgZFF_X2[12:12]),.O(Y_out_double_2_4_axb_12));
defparam Y_out_double_2_4_axb_12_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_13_cZ(.I0(Y_out_double_2_7[13:13]),.I1(pgZFF_X2[13:13]),.O(Y_out_double_2_4_axb_13));
defparam Y_out_double_2_4_axb_13_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_14_cZ(.I0(Y_out_double_2_7[14:14]),.I1(pgZFF_X2[14:14]),.O(Y_out_double_2_4_axb_14));
defparam Y_out_double_2_4_axb_14_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_15_cZ(.I0(Y_out_double_2_7[15:15]),.I1(pgZFF_X2[16:16]),.O(Y_out_double_2_4_axb_15));
defparam Y_out_double_2_4_axb_15_cZ.INIT=4'h6;
  LUT2 Y_out_double_2_4_axb_16_cZ(.I0(Y_out_double_2_7[17:17]),.I1(pgZFF_X2[16:16]),.O(Y_out_double_2_4_axb_16));
defparam Y_out_double_2_4_axb_16_cZ.INIT=4'h6;
  LUT2 un9_ac0_185(.I0(un9_8[6:6]),.I1(un9_10[8:8]),.O(un9_ac0_105));
defparam un9_ac0_185.INIT=4'h1;
  LUT2 un9_8_axb_29_cZ(.I0(ZFF_Y1[15:15]),.I1(ZFF_Y1[16:16]),.O(un9_8_axb_29));
defparam un9_8_axb_29_cZ.INIT=4'h9;
  LUT3 ZFF_Y1_8_rep1_RNI21EM(.I0(ZFF_Y1_5_rep1),.I1(ZFF_Y1_8_rep1),.I2(ZFF_Y1_fast[7:7]),.O(un9_6_0_axb_8));
defparam ZFF_Y1_8_rep1_RNI21EM.INIT=8'h36;
  LUT1 un6_0_6_cry_22_outextlut(.I0(GND),.O(un6_0_6_1[28:28]));
defparam un6_0_6_cry_22_outextlut.INIT=2'h3;
  LUT1 un9_6_0_cry_46_outextlut(.I0(GND),.O(un9_6_1[47:47]));
defparam un9_6_0_cry_46_outextlut.INIT=2'h3;
  LUT1 un9_8_cry_37_outextlut(.I0(GND),.O(un9_8_1[46:46]));
defparam un9_8_cry_37_outextlut.INIT=2'h3;
  LUT1 un9_10_cry_29_outextlut(.I0(GND),.O(un9_10_1[42:42]));
defparam un9_10_cry_29_outextlut.INIT=2'h3;
  LUT1 un10_6_cry_26_outextlut(.I0(GND),.O(un10_6_1[36:36]));
defparam un10_6_cry_26_outextlut.INIT=2'h3;
  LUT1 un8_0_6_cry_22_outextlut(.I0(GND),.O(un8_0_6_1[28:28]));
defparam un8_0_6_cry_22_outextlut.INIT=2'h3;
  LUT1 un7_0_6_cry_29_outextlut(.I0(GND),.O(un7_0_6_1[33:33]));
defparam un7_0_6_cry_29_outextlut.INIT=2'h3;
  LUT1 un7_0_8_cry_28_outextlut(.I0(GND),.O(un7_0_8_1[38:38]));
defparam un7_0_8_cry_28_outextlut.INIT=2'h3;
  LUT1 un6_0_8_cry_28_outextlut(.I0(GND),.O(un6_0_8_1[39:39]));
defparam un6_0_8_cry_28_outextlut.INIT=2'h3;
  LUT1 un8_0_8_cry_28_outextlut(.I0(GND),.O(un8_0_8_1[39:39]));
defparam un8_0_8_cry_28_outextlut.INIT=2'h3;
  LUT1 un6_0_9_cry_26_outextlut(.I0(GND),.O(un6_0_9_1[42:42]));
defparam un6_0_9_cry_26_outextlut.INIT=2'h3;
  LUT1 un8_0_9_cry_26_outextlut(.I0(GND),.O(un8_0_9_1[42:42]));
defparam un8_0_9_cry_26_outextlut.INIT=2'h3;
  LUT1 un9_11_cry_24_outextlut(.I0(GND),.O(un9_11_1[46:46]));
defparam un9_11_cry_24_outextlut.INIT=2'h3;
  LUT1 un9_8_cry_29_outextlut(.I0(GND),.O(un9_8_cry_29_1));
defparam un9_8_cry_29_outextlut.INIT=2'h3;
  LUT1 un9_6_0_cry_8_outextlut(.I0(GND),.O(un9_6_0_cry_8_1));
defparam un9_6_0_cry_8_outextlut.INIT=2'h3;
  INV n_reset_RNIG8S(.I(n_reset),.O(n_reset_i));
  p_O_FDE desc162(.Q(Y_out[0:0]),.D(Y_out_double[0:0]),.C(clk),.CE(trunc_out),.E(p_desc162_p_O_FDE));
  p_O_FDE desc163(.Q(Y_out[1:1]),.D(Y_out_double[1:1]),.C(clk),.CE(trunc_out),.E(p_desc163_p_O_FDE));
  p_O_FDE desc164(.Q(Y_out[2:2]),.D(Y_out_double[2:2]),.C(clk),.CE(trunc_out),.E(p_desc164_p_O_FDE));
  p_O_FDE desc165(.Q(Y_out[3:3]),.D(Y_out_double[3:3]),.C(clk),.CE(trunc_out),.E(p_desc165_p_O_FDE));
  p_O_FDE desc166(.Q(Y_out[4:4]),.D(Y_out_double[4:4]),.C(clk),.CE(trunc_out),.E(p_desc166_p_O_FDE));
  p_O_FDE desc167(.Q(Y_out[5:5]),.D(Y_out_double[5:5]),.C(clk),.CE(trunc_out),.E(p_desc167_p_O_FDE));
  p_O_FDE desc168(.Q(Y_out[6:6]),.D(Y_out_double[6:6]),.C(clk),.CE(trunc_out),.E(p_desc168_p_O_FDE));
  p_O_FDE desc169(.Q(Y_out[7:7]),.D(Y_out_double[7:7]),.C(clk),.CE(trunc_out),.E(p_desc169_p_O_FDE));
  p_O_FDE desc170(.Q(Y_out[8:8]),.D(Y_out_double[8:8]),.C(clk),.CE(trunc_out),.E(p_desc170_p_O_FDE));
  p_O_FDE desc171(.Q(Y_out[9:9]),.D(Y_out_double[9:9]),.C(clk),.CE(trunc_out),.E(p_desc171_p_O_FDE));
  p_O_FDE desc172(.Q(Y_out[10:10]),.D(Y_out_double[10:10]),.C(clk),.CE(trunc_out),.E(p_desc172_p_O_FDE));
  p_O_FDE desc173(.Q(Y_out[11:11]),.D(Y_out_double[11:11]),.C(clk),.CE(trunc_out),.E(p_desc173_p_O_FDE));
  p_O_FDE desc174(.Q(Y_out[12:12]),.D(Y_out_double[12:12]),.C(clk),.CE(trunc_out),.E(p_desc174_p_O_FDE));
  p_O_FDE desc175(.Q(Y_out[13:13]),.D(Y_out_double[13:13]),.C(clk),.CE(trunc_out),.E(p_desc175_p_O_FDE));
  p_O_FDE desc176(.Q(Y_out[14:14]),.D(Y_out_double[14:14]),.C(clk),.CE(trunc_out),.E(p_desc176_p_O_FDE));
  p_O_FDE desc177(.Q(Y_out[15:15]),.D(Y_out_double[15:15]),.C(clk),.CE(trunc_out),.E(p_desc177_p_O_FDE));
  p_O_FDE desc178(.Q(Y_out[16:16]),.D(Y_out_double[16:16]),.C(clk),.CE(trunc_out),.E(p_desc178_p_O_FDE));
  p_O_FDE desc179(.Q(Y_out[17:17]),.D(Y_out_double[17:17]),.C(clk),.CE(trunc_out),.E(p_desc179_p_O_FDE));
  p_O_FDCE desc180(.Q(un9_10[8:8]),.D(Y_out_double[0:0]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc180_p_O_FDCE));
  p_O_FDCE desc181(.Q(un9_8[6:6]),.D(Y_out_double[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc181_p_O_FDCE));
  p_O_FDCE desc182(.Q(un9_8[7:7]),.D(Y_out_double[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc182_p_O_FDCE));
  p_O_FDCE desc183(.Q(ZFF_Y1[3:3]),.D(Y_out_double[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc183_p_O_FDCE));
  p_O_FDCE desc184(.Q(ZFF_Y1[4:4]),.D(Y_out_double[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc184_p_O_FDCE));
  p_O_FDCE desc185(.Q(ZFF_Y1[5:5]),.D(Y_out_double[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc185_p_O_FDCE));
  p_O_FDCE desc186(.Q(ZFF_Y1[6:6]),.D(Y_out_double[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc186_p_O_FDCE));
  p_O_FDCE desc187(.Q(ZFF_Y1[7:7]),.D(Y_out_double[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc187_p_O_FDCE));
  p_O_FDCE desc188(.Q(ZFF_Y1[8:8]),.D(Y_out_double[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc188_p_O_FDCE));
  p_O_FDCE desc189(.Q(ZFF_Y1[9:9]),.D(Y_out_double[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc189_p_O_FDCE));
  p_O_FDCE desc190(.Q(un9_11[22:22]),.D(Y_out_double[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc190_p_O_FDCE));
  p_O_FDCE desc191(.Q(un9_11[23:23]),.D(Y_out_double[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc191_p_O_FDCE));
  p_O_FDCE desc192(.Q(un9_11[24:24]),.D(Y_out_double[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc192_p_O_FDCE));
  p_O_FDCE desc193(.Q(un9_11[25:25]),.D(Y_out_double[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc193_p_O_FDCE));
  p_O_FDCE desc194(.Q(un9_11[26:26]),.D(Y_out_double[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc194_p_O_FDCE));
  p_O_FDCE desc195(.Q(ZFF_Y1[15:15]),.D(Y_out_double[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc195_p_O_FDCE));
  p_O_FDCE desc196(.Q(ZFF_Y1[16:16]),.D(Y_out_double[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc196_p_O_FDCE));
  p_O_FDCE desc197(.Q(ZFF_Y1[17:17]),.D(Y_out_double[17:17]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc197_p_O_FDCE));
  p_O_FDE desc198(.Q(Y_out_double[0:0]),.D(Y_out_double_2[0:0]),.C(clk),.CE(sum_stg_a),.E(p_desc198_p_O_FDE));
  p_O_FDE desc199(.Q(Y_out_double[1:1]),.D(Y_out_double_2[1:1]),.C(clk),.CE(sum_stg_a),.E(p_desc199_p_O_FDE));
  p_O_FDE desc200(.Q(Y_out_double[2:2]),.D(Y_out_double_2[2:2]),.C(clk),.CE(sum_stg_a),.E(p_desc200_p_O_FDE));
  p_O_FDE desc201(.Q(Y_out_double[3:3]),.D(Y_out_double_2[3:3]),.C(clk),.CE(sum_stg_a),.E(p_desc201_p_O_FDE));
  p_O_FDE desc202(.Q(Y_out_double[4:4]),.D(Y_out_double_2[4:4]),.C(clk),.CE(sum_stg_a),.E(p_desc202_p_O_FDE));
  p_O_FDE desc203(.Q(Y_out_double[5:5]),.D(Y_out_double_2[5:5]),.C(clk),.CE(sum_stg_a),.E(p_desc203_p_O_FDE));
  p_O_FDE desc204(.Q(Y_out_double[6:6]),.D(Y_out_double_2[6:6]),.C(clk),.CE(sum_stg_a),.E(p_desc204_p_O_FDE));
  p_O_FDE desc205(.Q(Y_out_double[7:7]),.D(Y_out_double_2[7:7]),.C(clk),.CE(sum_stg_a),.E(p_desc205_p_O_FDE));
  p_O_FDE desc206(.Q(Y_out_double[8:8]),.D(Y_out_double_2[8:8]),.C(clk),.CE(sum_stg_a),.E(p_desc206_p_O_FDE));
  p_O_FDE desc207(.Q(Y_out_double[9:9]),.D(Y_out_double_2[9:9]),.C(clk),.CE(sum_stg_a),.E(p_desc207_p_O_FDE));
  p_O_FDE desc208(.Q(Y_out_double[10:10]),.D(Y_out_double_2[10:10]),.C(clk),.CE(sum_stg_a),.E(p_desc208_p_O_FDE));
  p_O_FDE desc209(.Q(Y_out_double[11:11]),.D(Y_out_double_2[11:11]),.C(clk),.CE(sum_stg_a),.E(p_desc209_p_O_FDE));
  p_O_FDE desc210(.Q(Y_out_double[12:12]),.D(Y_out_double_2[12:12]),.C(clk),.CE(sum_stg_a),.E(p_desc210_p_O_FDE));
  p_O_FDE desc211(.Q(Y_out_double[13:13]),.D(Y_out_double_2[13:13]),.C(clk),.CE(sum_stg_a),.E(p_desc211_p_O_FDE));
  p_O_FDE desc212(.Q(Y_out_double[14:14]),.D(Y_out_double_2[14:14]),.C(clk),.CE(sum_stg_a),.E(p_desc212_p_O_FDE));
  p_O_FDE desc213(.Q(Y_out_double[15:15]),.D(Y_out_double_2[15:15]),.C(clk),.CE(sum_stg_a),.E(p_desc213_p_O_FDE));
  p_O_FDE desc214(.Q(Y_out_double[16:16]),.D(Y_out_double_2[16:16]),.C(clk),.CE(sum_stg_a),.E(p_desc214_p_O_FDE));
  p_O_FDE desc215(.Q(Y_out_double[17:17]),.D(Y_out_double_2[17:17]),.C(clk),.CE(sum_stg_a),.E(p_desc215_p_O_FDE));
  p_O_FDE desc216(.Q(pgZFF_X1[0:0]),.D(pgZFF_X1_quad[30:30]),.C(clk),.CE(trunc_prods),.E(p_desc216_p_O_FDE));
  p_O_FDE desc217(.Q(pgZFF_X1[1:1]),.D(pgZFF_X1_quad[31:31]),.C(clk),.CE(trunc_prods),.E(p_desc217_p_O_FDE));
  p_O_FDE desc218(.Q(pgZFF_X1[2:2]),.D(pgZFF_X1_quad[32:32]),.C(clk),.CE(trunc_prods),.E(p_desc218_p_O_FDE));
  p_O_FDE desc219(.Q(pgZFF_X1[3:3]),.D(pgZFF_X1_quad[33:33]),.C(clk),.CE(trunc_prods),.E(p_desc219_p_O_FDE));
  p_O_FDE desc220(.Q(pgZFF_X1[4:4]),.D(pgZFF_X1_quad[34:34]),.C(clk),.CE(trunc_prods),.E(p_desc220_p_O_FDE));
  p_O_FDE desc221(.Q(pgZFF_X1[5:5]),.D(pgZFF_X1_quad[35:35]),.C(clk),.CE(trunc_prods),.E(p_desc221_p_O_FDE));
  p_O_FDE desc222(.Q(pgZFF_X1[6:6]),.D(pgZFF_X1_quad[36:36]),.C(clk),.CE(trunc_prods),.E(p_desc222_p_O_FDE));
  p_O_FDE desc223(.Q(pgZFF_X1[7:7]),.D(pgZFF_X1_quad[37:37]),.C(clk),.CE(trunc_prods),.E(p_desc223_p_O_FDE));
  p_O_FDE desc224(.Q(pgZFF_X1[8:8]),.D(pgZFF_X1_quad[38:38]),.C(clk),.CE(trunc_prods),.E(p_desc224_p_O_FDE));
  p_O_FDE desc225(.Q(pgZFF_X1[9:9]),.D(pgZFF_X1_quad[39:39]),.C(clk),.CE(trunc_prods),.E(p_desc225_p_O_FDE));
  p_O_FDE desc226(.Q(pgZFF_X1[10:10]),.D(pgZFF_X1_quad[40:40]),.C(clk),.CE(trunc_prods),.E(p_desc226_p_O_FDE));
  p_O_FDE desc227(.Q(pgZFF_X1[11:11]),.D(pgZFF_X1_quad[41:41]),.C(clk),.CE(trunc_prods),.E(p_desc227_p_O_FDE));
  p_O_FDE desc228(.Q(pgZFF_X1[12:12]),.D(pgZFF_X1_quad[42:42]),.C(clk),.CE(trunc_prods),.E(p_desc228_p_O_FDE));
  p_O_FDE desc229(.Q(pgZFF_X1[13:13]),.D(pgZFF_X1_quad[43:43]),.C(clk),.CE(trunc_prods),.E(p_desc229_p_O_FDE));
  p_O_FDE desc230(.Q(pgZFF_X1[14:14]),.D(pgZFF_X1_quad[44:44]),.C(clk),.CE(trunc_prods),.E(p_desc230_p_O_FDE));
  p_O_FDE desc231(.Q(pgZFF_X1[15:15]),.D(pgZFF_X1_quad[45:45]),.C(clk),.CE(trunc_prods),.E(p_desc231_p_O_FDE));
  p_O_FDE desc232(.Q(pgZFF_X1[17:17]),.D(pgZFF_X1_quad[47:47]),.C(clk),.CE(trunc_prods),.E(p_desc232_p_O_FDE));
  p_O_FDE desc233(.Q(pgZFF_X2[0:0]),.D(pgZFF_X2_quad[30:30]),.C(clk),.CE(trunc_prods),.E(p_desc233_p_O_FDE));
  p_O_FDE desc234(.Q(pgZFF_X2[1:1]),.D(pgZFF_X2_quad[31:31]),.C(clk),.CE(trunc_prods),.E(p_desc234_p_O_FDE));
  p_O_FDE desc235(.Q(pgZFF_X2[2:2]),.D(pgZFF_X2_quad[32:32]),.C(clk),.CE(trunc_prods),.E(p_desc235_p_O_FDE));
  p_O_FDE desc236(.Q(pgZFF_X2[3:3]),.D(pgZFF_X2_quad[33:33]),.C(clk),.CE(trunc_prods),.E(p_desc236_p_O_FDE));
  p_O_FDE desc237(.Q(pgZFF_X2[4:4]),.D(pgZFF_X2_quad[34:34]),.C(clk),.CE(trunc_prods),.E(p_desc237_p_O_FDE));
  p_O_FDE desc238(.Q(pgZFF_X2[5:5]),.D(pgZFF_X2_quad[35:35]),.C(clk),.CE(trunc_prods),.E(p_desc238_p_O_FDE));
  p_O_FDE desc239(.Q(pgZFF_X2[6:6]),.D(pgZFF_X2_quad[36:36]),.C(clk),.CE(trunc_prods),.E(p_desc239_p_O_FDE));
  p_O_FDE desc240(.Q(pgZFF_X2[7:7]),.D(pgZFF_X2_quad[37:37]),.C(clk),.CE(trunc_prods),.E(p_desc240_p_O_FDE));
  p_O_FDE desc241(.Q(pgZFF_X2[8:8]),.D(pgZFF_X2_quad[38:38]),.C(clk),.CE(trunc_prods),.E(p_desc241_p_O_FDE));
  p_O_FDE desc242(.Q(pgZFF_X2[9:9]),.D(pgZFF_X2_quad[39:39]),.C(clk),.CE(trunc_prods),.E(p_desc242_p_O_FDE));
  p_O_FDE desc243(.Q(pgZFF_X2[10:10]),.D(pgZFF_X2_quad[40:40]),.C(clk),.CE(trunc_prods),.E(p_desc243_p_O_FDE));
  p_O_FDE desc244(.Q(pgZFF_X2[11:11]),.D(pgZFF_X2_quad[41:41]),.C(clk),.CE(trunc_prods),.E(p_desc244_p_O_FDE));
  p_O_FDE desc245(.Q(pgZFF_X2[12:12]),.D(pgZFF_X2_quad[42:42]),.C(clk),.CE(trunc_prods),.E(p_desc245_p_O_FDE));
  p_O_FDE desc246(.Q(pgZFF_X2[13:13]),.D(pgZFF_X2_quad[43:43]),.C(clk),.CE(trunc_prods),.E(p_desc246_p_O_FDE));
  p_O_FDE desc247(.Q(pgZFF_X2[14:14]),.D(pgZFF_X2_quad[44:44]),.C(clk),.CE(trunc_prods),.E(p_desc247_p_O_FDE));
  p_O_FDE desc248(.Q(pgZFF_X2[16:16]),.D(pgZFF_X2_quad[46:46]),.C(clk),.CE(trunc_prods),.E(p_desc248_p_O_FDE));
  p_O_FDE desc249(.Q(pgZFF_X0[0:0]),.D(pgZFF_X0_quad[30:30]),.C(clk),.CE(trunc_prods),.E(p_desc249_p_O_FDE));
  p_O_FDE desc250(.Q(pgZFF_X0[1:1]),.D(pgZFF_X0_quad[31:31]),.C(clk),.CE(trunc_prods),.E(p_desc250_p_O_FDE));
  p_O_FDE desc251(.Q(pgZFF_X0[2:2]),.D(pgZFF_X0_quad[32:32]),.C(clk),.CE(trunc_prods),.E(p_desc251_p_O_FDE));
  p_O_FDE desc252(.Q(pgZFF_X0[3:3]),.D(pgZFF_X0_quad[33:33]),.C(clk),.CE(trunc_prods),.E(p_desc252_p_O_FDE));
  p_O_FDE desc253(.Q(pgZFF_X0[4:4]),.D(pgZFF_X0_quad[34:34]),.C(clk),.CE(trunc_prods),.E(p_desc253_p_O_FDE));
  p_O_FDE desc254(.Q(pgZFF_X0[5:5]),.D(pgZFF_X0_quad[35:35]),.C(clk),.CE(trunc_prods),.E(p_desc254_p_O_FDE));
  p_O_FDE desc255(.Q(pgZFF_X0[6:6]),.D(pgZFF_X0_quad[36:36]),.C(clk),.CE(trunc_prods),.E(p_desc255_p_O_FDE));
  p_O_FDE desc256(.Q(pgZFF_X0[7:7]),.D(pgZFF_X0_quad[37:37]),.C(clk),.CE(trunc_prods),.E(p_desc256_p_O_FDE));
  p_O_FDE desc257(.Q(pgZFF_X0[8:8]),.D(pgZFF_X0_quad[38:38]),.C(clk),.CE(trunc_prods),.E(p_desc257_p_O_FDE));
  p_O_FDE desc258(.Q(pgZFF_X0[9:9]),.D(pgZFF_X0_quad[39:39]),.C(clk),.CE(trunc_prods),.E(p_desc258_p_O_FDE));
  p_O_FDE desc259(.Q(pgZFF_X0[10:10]),.D(pgZFF_X0_quad[40:40]),.C(clk),.CE(trunc_prods),.E(p_desc259_p_O_FDE));
  p_O_FDE desc260(.Q(pgZFF_X0[11:11]),.D(pgZFF_X0_quad[41:41]),.C(clk),.CE(trunc_prods),.E(p_desc260_p_O_FDE));
  p_O_FDE desc261(.Q(pgZFF_X0[12:12]),.D(pgZFF_X0_quad[42:42]),.C(clk),.CE(trunc_prods),.E(p_desc261_p_O_FDE));
  p_O_FDE desc262(.Q(pgZFF_X0[13:13]),.D(pgZFF_X0_quad[43:43]),.C(clk),.CE(trunc_prods),.E(p_desc262_p_O_FDE));
  p_O_FDE desc263(.Q(pgZFF_X0[14:14]),.D(pgZFF_X0_quad[44:44]),.C(clk),.CE(trunc_prods),.E(p_desc263_p_O_FDE));
  p_O_FDE desc264(.Q(pgZFF_X0[16:16]),.D(pgZFF_X0_quad[46:46]),.C(clk),.CE(trunc_prods),.E(p_desc264_p_O_FDE));
  p_O_FDCE desc265(.Q(ZFF_X2[0:0]),.D(ZFF_X1[0:0]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc265_p_O_FDCE));
  p_O_FDCE desc266(.Q(ZFF_X2[1:1]),.D(ZFF_X1[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc266_p_O_FDCE));
  p_O_FDCE desc267(.Q(ZFF_X2[2:2]),.D(ZFF_X1[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc267_p_O_FDCE));
  p_O_FDCE desc268(.Q(ZFF_X2[3:3]),.D(ZFF_X1[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc268_p_O_FDCE));
  p_O_FDCE desc269(.Q(ZFF_X2[4:4]),.D(ZFF_X1[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc269_p_O_FDCE));
  p_O_FDCE desc270(.Q(ZFF_X2[5:5]),.D(ZFF_X1[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc270_p_O_FDCE));
  p_O_FDCE desc271(.Q(ZFF_X2[6:6]),.D(ZFF_X1[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc271_p_O_FDCE));
  p_O_FDCE desc272(.Q(ZFF_X2[7:7]),.D(ZFF_X1[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc272_p_O_FDCE));
  p_O_FDCE desc273(.Q(ZFF_X2[8:8]),.D(ZFF_X1[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc273_p_O_FDCE));
  p_O_FDCE desc274(.Q(ZFF_X2[9:9]),.D(ZFF_X1[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc274_p_O_FDCE));
  p_O_FDCE desc275(.Q(ZFF_X2[10:10]),.D(ZFF_X1[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc275_p_O_FDCE));
  p_O_FDCE desc276(.Q(ZFF_X2[11:11]),.D(ZFF_X1[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc276_p_O_FDCE));
  p_O_FDCE desc277(.Q(ZFF_X2[12:12]),.D(ZFF_X1[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc277_p_O_FDCE));
  p_O_FDCE desc278(.Q(ZFF_X2[13:13]),.D(ZFF_X1[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc278_p_O_FDCE));
  p_O_FDCE desc279(.Q(ZFF_X2[14:14]),.D(ZFF_X1[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc279_p_O_FDCE));
  p_O_FDCE desc280(.Q(ZFF_X2[15:15]),.D(ZFF_X1[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc280_p_O_FDCE));
  p_O_FDCE desc281(.Q(ZFF_X2[16:16]),.D(ZFF_X1[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc281_p_O_FDCE));
  p_O_FDCE desc282(.Q(ZFF_X1[0:0]),.D(ZFF_X0[0:0]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc282_p_O_FDCE));
  p_O_FDCE desc283(.Q(ZFF_X1[1:1]),.D(ZFF_X0[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc283_p_O_FDCE));
  p_O_FDCE desc284(.Q(ZFF_X1[2:2]),.D(ZFF_X0[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc284_p_O_FDCE));
  p_O_FDCE desc285(.Q(ZFF_X1[3:3]),.D(ZFF_X0[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc285_p_O_FDCE));
  p_O_FDCE desc286(.Q(ZFF_X1[4:4]),.D(ZFF_X0[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc286_p_O_FDCE));
  p_O_FDCE desc287(.Q(ZFF_X1[5:5]),.D(ZFF_X0[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc287_p_O_FDCE));
  p_O_FDCE desc288(.Q(ZFF_X1[6:6]),.D(ZFF_X0[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc288_p_O_FDCE));
  p_O_FDCE desc289(.Q(ZFF_X1[7:7]),.D(ZFF_X0[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc289_p_O_FDCE));
  p_O_FDCE desc290(.Q(ZFF_X1[8:8]),.D(ZFF_X0[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc290_p_O_FDCE));
  p_O_FDCE desc291(.Q(ZFF_X1[9:9]),.D(ZFF_X0[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc291_p_O_FDCE));
  p_O_FDCE desc292(.Q(ZFF_X1[10:10]),.D(ZFF_X0[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc292_p_O_FDCE));
  p_O_FDCE desc293(.Q(ZFF_X1[11:11]),.D(ZFF_X0[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc293_p_O_FDCE));
  p_O_FDCE desc294(.Q(ZFF_X1[12:12]),.D(ZFF_X0[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc294_p_O_FDCE));
  p_O_FDCE desc295(.Q(ZFF_X1[13:13]),.D(ZFF_X0[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc295_p_O_FDCE));
  p_O_FDCE desc296(.Q(ZFF_X1[14:14]),.D(ZFF_X0[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc296_p_O_FDCE));
  p_O_FDCE desc297(.Q(ZFF_X1[15:15]),.D(ZFF_X0[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc297_p_O_FDCE));
  p_O_FDCE desc298(.Q(ZFF_X1[16:16]),.D(ZFF_X0[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc298_p_O_FDCE));
  p_O_FDCE desc299(.Q(ZFF_Y2[0:0]),.D(un9_10[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc299_p_O_FDCE));
  p_O_FDCE desc300(.Q(ZFF_Y2[1:1]),.D(un9_8[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc300_p_O_FDCE));
  p_O_FDCE desc301(.Q(ZFF_Y2[2:2]),.D(un9_8[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc301_p_O_FDCE));
  p_O_FDCE desc302(.Q(ZFF_Y2[3:3]),.D(ZFF_Y1[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc302_p_O_FDCE));
  p_O_FDCE desc303(.Q(ZFF_Y2[4:4]),.D(ZFF_Y1[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc303_p_O_FDCE));
  p_O_FDCE desc304(.Q(ZFF_Y2[5:5]),.D(ZFF_Y1[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc304_p_O_FDCE));
  p_O_FDCE desc305(.Q(ZFF_Y2[6:6]),.D(ZFF_Y1[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc305_p_O_FDCE));
  p_O_FDCE desc306(.Q(ZFF_Y2[7:7]),.D(ZFF_Y1[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc306_p_O_FDCE));
  p_O_FDCE desc307(.Q(ZFF_Y2[8:8]),.D(ZFF_Y1[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc307_p_O_FDCE));
  p_O_FDCE desc308(.Q(ZFF_Y2[9:9]),.D(ZFF_Y1[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc308_p_O_FDCE));
  p_O_FDCE desc309(.Q(ZFF_Y2[10:10]),.D(un9_11[22:22]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc309_p_O_FDCE));
  p_O_FDCE desc310(.Q(ZFF_Y2[11:11]),.D(un9_11[23:23]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc310_p_O_FDCE));
  p_O_FDCE desc311(.Q(ZFF_Y2[12:12]),.D(un9_11[24:24]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc311_p_O_FDCE));
  p_O_FDCE desc312(.Q(ZFF_Y2[13:13]),.D(un9_11[25:25]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc312_p_O_FDCE));
  p_O_FDCE desc313(.Q(ZFF_Y2[14:14]),.D(un9_11[26:26]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc313_p_O_FDCE));
  p_O_FDCE desc314(.Q(ZFF_Y2[15:15]),.D(ZFF_Y1[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc314_p_O_FDCE));
  p_O_FDCE desc315(.Q(ZFF_Y2[16:16]),.D(ZFF_Y1[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc315_p_O_FDCE));
  p_O_FDCE desc316(.Q(ZFF_Y2[17:17]),.D(ZFF_Y1[17:17]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc316_p_O_FDCE));
  p_O_FDCE desc317(.Q(ZFF_X0[0:0]),.D(X_in[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc317_p_O_FDCE));
  p_O_FDCE desc318(.Q(ZFF_X0[1:1]),.D(X_in[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc318_p_O_FDCE));
  p_O_FDCE desc319(.Q(ZFF_X0[2:2]),.D(X_in[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc319_p_O_FDCE));
  p_O_FDCE desc320(.Q(ZFF_X0[3:3]),.D(X_in[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc320_p_O_FDCE));
  p_O_FDCE desc321(.Q(ZFF_X0[4:4]),.D(X_in[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc321_p_O_FDCE));
  p_O_FDCE desc322(.Q(ZFF_X0[5:5]),.D(X_in[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc322_p_O_FDCE));
  p_O_FDCE desc323(.Q(ZFF_X0[6:6]),.D(X_in[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc323_p_O_FDCE));
  p_O_FDCE desc324(.Q(ZFF_X0[7:7]),.D(X_in[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc324_p_O_FDCE));
  p_O_FDCE desc325(.Q(ZFF_X0[8:8]),.D(X_in[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc325_p_O_FDCE));
  p_O_FDCE desc326(.Q(ZFF_X0[9:9]),.D(X_in[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc326_p_O_FDCE));
  p_O_FDCE desc327(.Q(ZFF_X0[10:10]),.D(X_in[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc327_p_O_FDCE));
  p_O_FDCE desc328(.Q(ZFF_X0[11:11]),.D(X_in[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc328_p_O_FDCE));
  p_O_FDCE desc329(.Q(ZFF_X0[12:12]),.D(X_in[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc329_p_O_FDCE));
  p_O_FDCE desc330(.Q(ZFF_X0[13:13]),.D(X_in[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc330_p_O_FDCE));
  p_O_FDCE desc331(.Q(ZFF_X0[14:14]),.D(X_in[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc331_p_O_FDCE));
  p_O_FDCE desc332(.Q(ZFF_X0[15:15]),.D(X_in[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc332_p_O_FDCE));
  p_O_FDCE desc333(.Q(ZFF_X0[16:16]),.D(X_in[17:17]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc333_p_O_FDCE));
  p_O_FDC desc334(.Q(q_reg[2:2]),.D(q_next[2:2]),.C(clk),.CLR(n_reset_i),.E(p_desc334_p_O_FDC));
  p_O_FDC desc335(.Q(q_reg[1:1]),.D(q_next[1:1]),.C(clk),.CLR(n_reset_i),.E(p_desc335_p_O_FDC));
  p_O_FDC desc336(.Q(q_reg[0:0]),.D(q_next[0:0]),.C(clk),.CLR(n_reset_i),.E(p_desc336_p_O_FDC));
  p_O_FDC desc337(.Q(state_reg),.D(state_next),.C(clk),.CLR(n_reset_i),.E(p_desc337_p_O_FDC));
  p_O_FDP state_reg_ret_Z(.Q(q_reg_i_1[2:2]),.D(q_next_i[2:2]),.C(clk),.PRE(n_reset_i),.E(p_state_reg_ret_Z_p_O_FDP));
  p_O_FDP state_reg_ret_1_Z(.Q(q_reg_i_1[1:1]),.D(q_next_i[1:1]),.C(clk),.PRE(n_reset_i),.E(p_state_reg_ret_1_Z_p_O_FDP));
  p_O_FDP state_reg_ret_2_Z(.Q(q_reg_i_1[0:0]),.D(q_next_i[0:0]),.C(clk),.PRE(n_reset_i),.E(p_state_reg_ret_2_Z_p_O_FDP));
  p_O_FDP state_reg_ret_4_Z(.Q(state_reg_ret_4),.D(un7_q_reg_reti),.C(clk),.PRE(n_reset_i),.E(p_state_reg_ret_4_Z_p_O_FDP));
  p_O_FDC state_reg_ret_5_Z(.Q(un1_q_reg_2_c),.D(un1_q_reg_2_reti),.C(clk),.CLR(n_reset_i),.E(p_state_reg_ret_5_Z_p_O_FDC));
  p_O_FDCE desc338(.Q(un9_10_fast[8:8]),.D(Y_out_double[0:0]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc338_p_O_FDCE));
  p_O_FDCE ZFF_Y1_0_rep1_Z(.Q(un9_10_8_rep1),.D(Y_out_double[0:0]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_0_rep1_Z_p_O_FDCE));
  p_O_FDCE desc339(.Q(ZFF_Y1_fast[15:15]),.D(Y_out_double[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc339_p_O_FDCE));
  p_O_FDCE ZFF_Y1_15_rep1_Z(.Q(ZFF_Y1_15_rep1),.D(Y_out_double[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_15_rep1_Z_p_O_FDCE));
  p_O_FDCE desc340(.Q(ZFF_X0_fast[7:7]),.D(X_in[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc340_p_O_FDCE));
  p_O_FDCE ZFF_X0_7_rep1_Z(.Q(ZFF_X0_7_rep1),.D(X_in[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_7_rep1_Z_p_O_FDCE));
  p_O_FDCE desc341(.Q(ZFF_X0_fast[8:8]),.D(X_in[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc341_p_O_FDCE));
  p_O_FDCE desc342(.Q(ZFF_X2_fast[8:8]),.D(ZFF_X1[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc342_p_O_FDCE));
  p_O_FDCE desc343(.Q(ZFF_X2_fast[7:7]),.D(ZFF_X1[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc343_p_O_FDCE));
  p_O_FDCE desc344(.Q(ZFF_Y1_fast[16:16]),.D(Y_out_double[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc344_p_O_FDCE));
  p_O_FDCE ZFF_Y1_16_rep1_Z(.Q(ZFF_Y1_16_rep1),.D(Y_out_double[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_16_rep1_Z_p_O_FDCE));
  p_O_FDCE desc345(.Q(ZFF_X0_fast[6:6]),.D(X_in[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc345_p_O_FDCE));
  p_O_FDCE ZFF_X0_6_rep1_Z(.Q(ZFF_X0_6_rep1),.D(X_in[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_6_rep1_Z_p_O_FDCE));
  p_O_FDCE desc346(.Q(ZFF_X0_fast[5:5]),.D(X_in[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc346_p_O_FDCE));
  p_O_FDCE desc347(.Q(un9_8_fast[7:7]),.D(Y_out_double[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc347_p_O_FDCE));
  p_O_FDCE ZFF_Y1_2_rep1_Z(.Q(un9_8_7_rep1),.D(Y_out_double[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_2_rep1_Z_p_O_FDCE));
  p_O_FDCE desc348(.Q(ZFF_X2_fast[5:5]),.D(ZFF_X1[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc348_p_O_FDCE));
  p_O_FDCE desc349(.Q(ZFF_X0_fast[10:10]),.D(X_in[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc349_p_O_FDCE));
  p_O_FDCE ZFF_X0_10_rep1_Z(.Q(ZFF_X0_10_rep1),.D(X_in[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_10_rep1_Z_p_O_FDCE));
  p_O_FDCE desc350(.Q(ZFF_X0_fast[11:11]),.D(X_in[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc350_p_O_FDCE));
  p_O_FDCE ZFF_X0_11_rep1_Z(.Q(ZFF_X0_11_rep1),.D(X_in[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_11_rep1_Z_p_O_FDCE));
  p_O_FDCE desc351(.Q(ZFF_X0_fast[12:12]),.D(X_in[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc351_p_O_FDCE));
  p_O_FDCE ZFF_X0_12_rep1_Z(.Q(ZFF_X0_12_rep1),.D(X_in[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_12_rep1_Z_p_O_FDCE));
  p_O_FDCE desc352(.Q(ZFF_X2_fast[6:6]),.D(ZFF_X1[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc352_p_O_FDCE));
  p_O_FDCE ZFF_X2_6_rep1_Z(.Q(ZFF_X2_6_rep1),.D(ZFF_X1[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X2_6_rep1_Z_p_O_FDCE));
  p_O_FDCE desc353(.Q(ZFF_X0_fast[4:4]),.D(X_in[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc353_p_O_FDCE));
  p_O_FDCE ZFF_X0_4_rep1_Z(.Q(ZFF_X0_4_rep1),.D(X_in[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_4_rep1_Z_p_O_FDCE));
  p_O_FDCE desc354(.Q(ZFF_X2_fast[11:11]),.D(ZFF_X1[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc354_p_O_FDCE));
  p_O_FDCE desc355(.Q(ZFF_X2_fast[12:12]),.D(ZFF_X1[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc355_p_O_FDCE));
  p_O_FDCE desc356(.Q(ZFF_X0_fast[9:9]),.D(X_in[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc356_p_O_FDCE));
  p_O_FDCE desc357(.Q(ZFF_X2_fast[10:10]),.D(ZFF_X1[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc357_p_O_FDCE));
  p_O_FDCE ZFF_X2_10_rep1_Z(.Q(ZFF_X2_10_rep1),.D(ZFF_X1[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X2_10_rep1_Z_p_O_FDCE));
  p_O_FDCE desc358(.Q(ZFF_X0_fast[2:2]),.D(X_in[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc358_p_O_FDCE));
  p_O_FDCE ZFF_X0_2_rep1_Z(.Q(ZFF_X0_2_rep1),.D(X_in[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_2_rep1_Z_p_O_FDCE));
  p_O_FDCE desc359(.Q(ZFF_X0_fast[1:1]),.D(X_in[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc359_p_O_FDCE));
  p_O_FDCE ZFF_X0_1_rep1_Z(.Q(ZFF_X0_1_rep1),.D(X_in[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_1_rep1_Z_p_O_FDCE));
  p_O_FDCE desc360(.Q(un9_8_fast[6:6]),.D(Y_out_double[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc360_p_O_FDCE));
  p_O_FDCE ZFF_Y1_1_rep1_Z(.Q(un9_8_6_rep1),.D(Y_out_double[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_1_rep1_Z_p_O_FDCE));
  p_O_FDCE desc361(.Q(ZFF_X2_fast[4:4]),.D(ZFF_X1[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc361_p_O_FDCE));
  p_O_FDCE desc362(.Q(ZFF_X2_fast[9:9]),.D(ZFF_X1[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc362_p_O_FDCE));
  p_O_FDCE desc363(.Q(ZFF_X2_fast[1:1]),.D(ZFF_X1[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc363_p_O_FDCE));
  p_O_FDCE desc364(.Q(ZFF_X2_fast[2:2]),.D(ZFF_X1[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc364_p_O_FDCE));
  p_O_FDCE ZFF_X2_2_rep1_Z(.Q(ZFF_X2_2_rep1),.D(ZFF_X1[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X2_2_rep1_Z_p_O_FDCE));
  p_O_FDCE desc365(.Q(ZFF_X0_fast[3:3]),.D(X_in[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc365_p_O_FDCE));
  p_O_FDCE ZFF_X0_3_rep1_Z(.Q(ZFF_X0_3_rep1),.D(X_in[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_3_rep1_Z_p_O_FDCE));
  p_O_FDCE desc366(.Q(ZFF_X0_fast[13:13]),.D(X_in[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc366_p_O_FDCE));
  p_O_FDCE desc367(.Q(ZFF_X2_fast[3:3]),.D(ZFF_X1[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc367_p_O_FDCE));
  p_O_FDCE ZFF_X2_3_rep1_Z(.Q(ZFF_X2_3_rep1),.D(ZFF_X1[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X2_3_rep1_Z_p_O_FDCE));
  p_O_FDCE desc368(.Q(ZFF_Y1_fast[4:4]),.D(Y_out_double[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc368_p_O_FDCE));
  p_O_FDCE ZFF_Y1_4_rep1_Z(.Q(ZFF_Y1_4_rep1),.D(Y_out_double[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_4_rep1_Z_p_O_FDCE));
  p_O_FDCE desc369(.Q(ZFF_X2_fast[13:13]),.D(ZFF_X1[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc369_p_O_FDCE));
  p_O_FDCE desc370(.Q(ZFF_Y1_fast[3:3]),.D(Y_out_double[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc370_p_O_FDCE));
  p_O_FDCE ZFF_Y1_3_rep1_Z(.Q(ZFF_Y1_3_rep1),.D(Y_out_double[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_3_rep1_Z_p_O_FDCE));
  p_O_FDCE desc371(.Q(ZFF_X0_fast[0:0]),.D(X_in[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc371_p_O_FDCE));
  p_O_FDCE desc372(.Q(ZFF_X2_fast[0:0]),.D(ZFF_X1[0:0]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc372_p_O_FDCE));
  p_O_FDCE desc373(.Q(ZFF_Y1_fast[5:5]),.D(Y_out_double[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc373_p_O_FDCE));
  p_O_FDCE ZFF_Y1_5_rep1_Z(.Q(ZFF_Y1_5_rep1),.D(Y_out_double[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_5_rep1_Z_p_O_FDCE));
  p_O_FDCE desc374(.Q(ZFF_X2_fast[14:14]),.D(ZFF_X1[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc374_p_O_FDCE));
  p_O_FDCE ZFF_X2_14_rep1_Z(.Q(ZFF_X2_14_rep1),.D(ZFF_X1[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X2_14_rep1_Z_p_O_FDCE));
  p_O_FDCE desc375(.Q(ZFF_X0_fast[14:14]),.D(X_in[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc375_p_O_FDCE));
  p_O_FDCE ZFF_X0_14_rep1_Z(.Q(ZFF_X0_14_rep1),.D(X_in[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_14_rep1_Z_p_O_FDCE));
  p_O_FDCE desc376(.Q(ZFF_X0_fast[15:15]),.D(X_in[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc376_p_O_FDCE));
  p_O_FDCE ZFF_X0_15_rep1_Z(.Q(ZFF_X0_15_rep1),.D(X_in[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_15_rep1_Z_p_O_FDCE));
  p_O_FDCE desc377(.Q(ZFF_X2_fast[15:15]),.D(ZFF_X1[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc377_p_O_FDCE));
  p_O_FDCE ZFF_X2_15_rep1_Z(.Q(ZFF_X2_15_rep1),.D(ZFF_X1[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X2_15_rep1_Z_p_O_FDCE));
  p_O_FDCE desc378(.Q(ZFF_Y1_fast[6:6]),.D(Y_out_double[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc378_p_O_FDCE));
  p_O_FDCE ZFF_Y1_6_rep1_Z(.Q(ZFF_Y1_6_rep1),.D(Y_out_double[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_6_rep1_Z_p_O_FDCE));
  p_O_FDCE desc379(.Q(un9_11_fast[25:25]),.D(Y_out_double[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc379_p_O_FDCE));
  p_O_FDCE ZFF_Y1_13_rep1_Z(.Q(un9_11_25_rep1),.D(Y_out_double[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_13_rep1_Z_p_O_FDCE));
  p_O_FDCE desc380(.Q(ZFF_Y1_fast[7:7]),.D(Y_out_double[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc380_p_O_FDCE));
  p_O_FDCE ZFF_Y1_7_rep1_Z(.Q(ZFF_Y1_7_rep1),.D(Y_out_double[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_7_rep1_Z_p_O_FDCE));
  p_O_FDCE desc381(.Q(un9_11_fast[26:26]),.D(Y_out_double[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc381_p_O_FDCE));
  p_O_FDCE ZFF_Y1_14_rep1_Z(.Q(un9_11_26_rep1),.D(Y_out_double[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_14_rep1_Z_p_O_FDCE));
  p_O_FDCE desc382(.Q(ZFF_X1_fast[3:3]),.D(ZFF_X0[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc382_p_O_FDCE));
  p_O_FDCE ZFF_X1_3_rep1_Z(.Q(ZFF_X1_3_rep1),.D(ZFF_X0[3:3]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_3_rep1_Z_p_O_FDCE));
  p_O_FDCE desc383(.Q(ZFF_X1_fast[0:0]),.D(ZFF_X0[0:0]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc383_p_O_FDCE));
  p_O_FDCE ZFF_X1_0_rep1_Z(.Q(ZFF_X1_0_rep1),.D(ZFF_X0[0:0]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_0_rep1_Z_p_O_FDCE));
  p_O_FDCE desc384(.Q(ZFF_Y1_fast[9:9]),.D(Y_out_double[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc384_p_O_FDCE));
  p_O_FDCE ZFF_Y1_9_rep1_Z(.Q(ZFF_Y1_9_rep1),.D(Y_out_double[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_9_rep1_Z_p_O_FDCE));
  p_O_FDCE desc385(.Q(ZFF_X1_fast[7:7]),.D(ZFF_X0[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc385_p_O_FDCE));
  p_O_FDCE ZFF_X1_7_rep1_Z(.Q(ZFF_X1_7_rep1),.D(ZFF_X0[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_7_rep1_Z_p_O_FDCE));
  p_O_FDCE desc386(.Q(ZFF_X1_fast[4:4]),.D(ZFF_X0[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc386_p_O_FDCE));
  p_O_FDCE ZFF_X1_4_rep1_Z(.Q(ZFF_X1_4_rep1),.D(ZFF_X0[4:4]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_4_rep1_Z_p_O_FDCE));
  p_O_FDCE desc387(.Q(ZFF_X1_fast[1:1]),.D(ZFF_X0[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc387_p_O_FDCE));
  p_O_FDCE ZFF_X1_1_rep1_Z(.Q(ZFF_X1_1_rep1),.D(ZFF_X0[1:1]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_1_rep1_Z_p_O_FDCE));
  p_O_FDCE desc388(.Q(un9_11_fast[22:22]),.D(Y_out_double[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc388_p_O_FDCE));
  p_O_FDCE ZFF_Y1_10_rep1_Z(.Q(un9_11_22_rep1),.D(Y_out_double[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_10_rep1_Z_p_O_FDCE));
  p_O_FDCE desc389(.Q(ZFF_X1_fast[8:8]),.D(ZFF_X0[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc389_p_O_FDCE));
  p_O_FDCE ZFF_X1_8_rep1_Z(.Q(ZFF_X1_8_rep1),.D(ZFF_X0[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_8_rep1_Z_p_O_FDCE));
  p_O_FDCE desc390(.Q(ZFF_X1_fast[9:9]),.D(ZFF_X0[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc390_p_O_FDCE));
  p_O_FDCE ZFF_X1_9_rep1_Z(.Q(ZFF_X1_9_rep1),.D(ZFF_X0[9:9]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_9_rep1_Z_p_O_FDCE));
  p_O_FDCE desc391(.Q(ZFF_X1_fast[11:11]),.D(ZFF_X0[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc391_p_O_FDCE));
  p_O_FDCE ZFF_X1_11_rep1_Z(.Q(ZFF_X1_11_rep1),.D(ZFF_X0[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_11_rep1_Z_p_O_FDCE));
  p_O_FDCE desc392(.Q(ZFF_X1_fast[15:15]),.D(ZFF_X0[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc392_p_O_FDCE));
  p_O_FDCE ZFF_X1_15_rep1_Z(.Q(ZFF_X1_15_rep1),.D(ZFF_X0[15:15]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_15_rep1_Z_p_O_FDCE));
  p_O_FDCE desc393(.Q(ZFF_X1_fast[2:2]),.D(ZFF_X0[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc393_p_O_FDCE));
  p_O_FDCE ZFF_X1_2_rep1_Z(.Q(ZFF_X1_2_rep1),.D(ZFF_X0[2:2]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_2_rep1_Z_p_O_FDCE));
  p_O_FDCE desc394(.Q(un9_11_fast[24:24]),.D(Y_out_double[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc394_p_O_FDCE));
  p_O_FDCE ZFF_Y1_12_rep1_Z(.Q(un9_11_24_rep1),.D(Y_out_double[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_12_rep1_Z_p_O_FDCE));
  p_O_FDCE desc395(.Q(ZFF_X0_fast[16:16]),.D(X_in[17:17]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc395_p_O_FDCE));
  p_O_FDCE ZFF_X0_16_rep1_Z(.Q(ZFF_X0_16_rep1),.D(X_in[17:17]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X0_16_rep1_Z_p_O_FDCE));
  p_O_FDCE desc396(.Q(ZFF_X2_fast[16:16]),.D(ZFF_X1[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc396_p_O_FDCE));
  p_O_FDCE desc397(.Q(ZFF_Y1_fast[17:17]),.D(Y_out_double[17:17]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc397_p_O_FDCE));
  p_O_FDCE ZFF_Y1_17_rep1_Z(.Q(ZFF_Y1_17_rep1),.D(Y_out_double[17:17]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_17_rep1_Z_p_O_FDCE));
  p_O_FDCE desc398(.Q(ZFF_X1_fast[5:5]),.D(ZFF_X0[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc398_p_O_FDCE));
  p_O_FDCE ZFF_X1_5_rep1_Z(.Q(ZFF_X1_5_rep1),.D(ZFF_X0[5:5]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_5_rep1_Z_p_O_FDCE));
  p_O_FDCE desc399(.Q(ZFF_Y1_fast[8:8]),.D(Y_out_double[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc399_p_O_FDCE));
  p_O_FDCE ZFF_Y1_8_rep1_Z(.Q(ZFF_Y1_8_rep1),.D(Y_out_double[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_8_rep1_Z_p_O_FDCE));
  p_O_FDCE desc400(.Q(ZFF_X1_fast[14:14]),.D(ZFF_X0[14:14]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc400_p_O_FDCE));
  p_O_FDCE desc401(.Q(ZFF_X1_fast[16:16]),.D(ZFF_X0[16:16]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc401_p_O_FDCE));
  p_O_FDCE desc402(.Q(ZFF_X1_fast[6:6]),.D(ZFF_X0[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc402_p_O_FDCE));
  p_O_FDCE ZFF_X1_6_rep1_Z(.Q(ZFF_X1_6_rep1),.D(ZFF_X0[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_6_rep1_Z_p_O_FDCE));
  p_O_FDCE desc403(.Q(ZFF_X1_fast[12:12]),.D(ZFF_X0[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc403_p_O_FDCE));
  p_O_FDCE ZFF_X1_12_rep1_Z(.Q(ZFF_X1_12_rep1),.D(ZFF_X0[12:12]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_12_rep1_Z_p_O_FDCE));
  p_O_FDCE desc404(.Q(ZFF_X1_fast[10:10]),.D(ZFF_X0[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc404_p_O_FDCE));
  p_O_FDCE ZFF_X1_10_rep1_Z(.Q(ZFF_X1_10_rep1),.D(ZFF_X0[10:10]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_10_rep1_Z_p_O_FDCE));
  p_O_FDCE desc405(.Q(ZFF_X1_fast[13:13]),.D(ZFF_X0[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc405_p_O_FDCE));
  p_O_FDCE ZFF_X1_13_rep1_Z(.Q(ZFF_X1_13_rep1),.D(ZFF_X0[13:13]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_X1_13_rep1_Z_p_O_FDCE));
  p_O_FDCE desc406(.Q(un9_11_fast[23:23]),.D(Y_out_double[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc406_p_O_FDCE));
  p_O_FDCE ZFF_Y1_11_rep1_Z(.Q(un9_11_23_rep1),.D(Y_out_double[11:11]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y1_11_rep1_Z_p_O_FDCE));
  p_O_FDCE desc407(.Q(ZFF_Y2_fast[8:8]),.D(ZFF_Y1[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc407_p_O_FDCE));
  p_O_FDCE ZFF_Y2_8_rep1_Z(.Q(ZFF_Y2_8_rep1),.D(ZFF_Y1[8:8]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y2_8_rep1_Z_p_O_FDCE));
  p_O_FDCE desc408(.Q(ZFF_Y2_fast[17:17]),.D(ZFF_Y1[17:17]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc408_p_O_FDCE));
  p_O_FDCE desc409(.Q(ZFF_Y2_fast[6:6]),.D(ZFF_Y1[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc409_p_O_FDCE));
  p_O_FDCE ZFF_Y2_6_rep1_Z(.Q(ZFF_Y2_6_rep1),.D(ZFF_Y1[6:6]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y2_6_rep1_Z_p_O_FDCE));
  p_O_FDCE desc410(.Q(ZFF_Y2_fast[7:7]),.D(ZFF_Y1[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc410_p_O_FDCE));
  p_O_FDCE ZFF_Y2_7_rep1_Z(.Q(ZFF_Y2_7_rep1),.D(ZFF_Y1[7:7]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y2_7_rep1_Z_p_O_FDCE));
  p_O_FDCE desc411(.Q(ZFF_Y2_fast[14:14]),.D(un9_11[26:26]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_desc411_p_O_FDCE));
  p_O_FDCE ZFF_Y2_14_rep1_Z(.Q(ZFF_Y2_14_rep1),.D(un9_11[26:26]),.C(clk),.CLR(n_reset_i),.CE(sample_trig),.E(p_ZFF_Y2_14_rep1_Z_p_O_FDCE));
  MUXCY_L un9_6_0_cry_8_outext(.DI(GND),.CI(un9_6_0_cry_8_0),.S(un9_6_0_cry_8_1),.LO(un9_6_0_cry_8));
  MUXCY_L un9_8_cry_29_outext(.DI(GND),.CI(un9_8_cry_29_0),.S(un9_8_cry_29_1),.LO(un9_8_cry_29));
  MUXCY un9_11_cry_24_outext(.DI(GND),.CI(un9_11_0[46:46]),.S(un9_11_1[46:46]),.O(un9_11[46:46]));
  MUXCY un8_0_9_cry_26_outext(.DI(GND),.CI(un8_0_9_0[42:42]),.S(un8_0_9_1[42:42]),.O(un8_0_9[42:42]));
  MUXCY un6_0_9_cry_26_outext(.DI(GND),.CI(un6_0_9_0[42:42]),.S(un6_0_9_1[42:42]),.O(un6_0_9[42:42]));
  MUXCY un8_0_8_cry_28_outext(.DI(GND),.CI(un8_0_8[38:38]),.S(un8_0_8_1[39:39]),.O(un8_0_8[39:39]));
  MUXCY un6_0_8_cry_28_outext(.DI(GND),.CI(un6_0_8[38:38]),.S(un6_0_8_1[39:39]),.O(un6_0_8[39:39]));
  MUXCY un7_0_8_cry_28_outext(.DI(GND),.CI(un7_0_8_0[38:38]),.S(un7_0_8_1[38:38]),.O(un7_0_8[38:38]));
  MUXCY un7_0_6_cry_29_outext(.DI(GND),.CI(un7_0_6_0[33:33]),.S(un7_0_6_1[33:33]),.O(un7_0_6[33:33]));
  MUXCY un8_0_6_cry_22_outext(.DI(GND),.CI(un8_0_6_0[28:28]),.S(un8_0_6_1[28:28]),.O(un8_0_6[28:28]));
  MUXCY un10_6_cry_26_outext(.DI(GND),.CI(un10_6_0[36:36]),.S(un10_6_1[36:36]),.O(un10_6[36:36]));
  MUXCY un9_10_cry_29_outext(.DI(GND),.CI(un9_10_0[42:42]),.S(un9_10_1[42:42]),.O(un9_10[42:42]));
  MUXCY un9_8_cry_37_outext(.DI(GND),.CI(un9_8[45:45]),.S(un9_8_1[46:46]),.O(un9_8[46:46]));
  MUXCY un9_6_0_cry_46_outext(.DI(GND),.CI(un9_6_0[47:47]),.S(un9_6_1[47:47]),.O(un9_6[47:47]));
  MUXCY un6_0_6_cry_22_outext(.DI(GND),.CI(un6_0_6_0[28:28]),.S(un6_0_6_1[28:28]),.O(un6_0_6[28:28]));
  MUXCY un9_6_0_cry_8_cZ(.DI(un9_6_0_cry_8_RNO),.CI(un9_6_0_cry_7),.S(un9_6_0_axb_8),.O(un9_6_0_cry_8_0));
  MUXCY un9_8_cry_29_cZ(.DI(ZFF_Y1[15:15]),.CI(un9_8_cry_28),.S(un9_8_axb_29),.O(un9_8_cry_29_0));
  LUT2_L un6_0_0_axb_42_N_2L1_cZ(.I0(un6_0_9[39:39]),.I1(un6_0_9[40:40]),.LO(un6_0_0_axb_42_N_2L1));
defparam un6_0_0_axb_42_N_2L1_cZ.INIT=4'h7;
  LUT6 un6_0_0_axb_42_cZ(.I0(ZFF_X0[16:16]),.I1(un6_0_9[42:42]),.I2(un6_0_9[41:41]),.I3(un6_0_9[38:38]),.I4(un6_0_8[38:38]),.I5(un6_0_0_axb_42_N_2L1),.O(un6_0_0_axb_42));
defparam un6_0_0_axb_42_cZ.INIT=64'h6969696963696663;
  LUT2_L un8_0_0_axb_42_N_2L1_cZ(.I0(un8_0_9[39:39]),.I1(un8_0_9[40:40]),.LO(un8_0_0_axb_42_N_2L1));
defparam un8_0_0_axb_42_N_2L1_cZ.INIT=4'h7;
  LUT6 un8_0_0_axb_42_cZ(.I0(ZFF_X2[16:16]),.I1(un8_0_9[42:42]),.I2(un8_0_9[41:41]),.I3(un8_0_9[38:38]),.I4(un8_0_8[38:38]),.I5(un8_0_0_axb_42_N_2L1),.O(un8_0_0_axb_42));
defparam un8_0_0_axb_42_cZ.INIT=64'h6969696963696663;
  LUT5 un10_axb_9_cZ(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[6:6]),.I2(ZFF_Y2[14:14]),.I3(ZFF_Y2[9:9]),.I4(un10_6[15:15]),.O(un10_axb_9));
defparam un10_axb_9_cZ.INIT=32'h59A6A659;
  LUT2 un10_19_cZ(.I0(ZFF_Y2_6_rep1),.I1(ZFF_Y2_14_rep1),.O(un10_19));
defparam un10_19_cZ.INIT=4'h9;
  LUT6 un9_cry_7_RNO_0(.I0(ZFF_Y1[7:7]),.I1(ZFF_Y1[6:6]),.I2(ZFF_Y1[3:3]),.I3(un9_10[8:8]),.I4(un9_8[9:9]),.I5(un9_6[9:9]),.O(un9_axb_7));
defparam un9_cry_7_RNO_0.INIT=64'h965569AA69AA9655;
  LUT5 un10_8_axb_23_cZ(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2[12:12]),.I2(ZFF_Y2[13:13]),.I3(ZFF_Y2[15:15]),.I4(ZFF_Y2[17:17]),.O(un10_8_axb_23));
defparam un10_8_axb_23_cZ.INIT=32'h87781EE1;
  LUT5 un10_8_axb_24_cZ(.I0(ZFF_Y2[14:14]),.I1(ZFF_Y2[13:13]),.I2(ZFF_Y2[16:16]),.I3(ZFF_Y2[15:15]),.I4(ZFF_Y2[17:17]),.O(un10_8_axb_24));
defparam un10_8_axb_24_cZ.INIT=32'h965A5A69;
  LUT4 un9_o5_7_cZ(.I0(ZFF_Y1[9:9]),.I1(ZFF_Y1[7:7]),.I2(un9_8[9:9]),.I3(un9_6_0_cry_8),.O(un9_o5_7));
defparam un9_o5_7_cZ.INIT=16'hB271;
  LUT5 un6_0_8_axb_11_cZ(.I0(ZFF_X0_fast[15:15]),.I1(ZFF_X0_fast[6:6]),.I2(ZFF_X0_fast[0:0]),.I3(ZFF_X0_1_rep1),.I4(ZFF_X0_fast[5:5]),.O(un6_0_8_axb_11));
defparam un6_0_8_axb_11_cZ.INIT=32'h936CC936;
  LUT6 desc412(.I0(ZFF_X0_fast[14:14]),.I1(ZFF_X0_fast[12:12]),.I2(ZFF_X0_fast[4:4]),.I3(ZFF_X0_fast[11:11]),.I4(ZFF_X0_fast[3:3]),.I5(ZFF_X0_fast[13:13]),.O(un6_0_8_axb_9));
defparam desc412.INIT=64'h9669969669699669;
  LUT6 desc413(.I0(ZFF_X0_fast[1:1]),.I1(ZFF_X0_fast[2:2]),.I2(ZFF_X0_fast[10:10]),.I3(ZFF_X0_fast[12:12]),.I4(ZFF_X0_fast[11:11]),.I5(ZFF_X0_fast[9:9]),.O(un6_0_8_axb_7));
defparam desc413.INIT=64'hC33C699669963CC3;
  LUT6 desc414(.I0(ZFF_X2_fast[14:14]),.I1(ZFF_X2_fast[15:15]),.I2(ZFF_X2_fast[0:0]),.I3(ZFF_X2_fast[4:4]),.I4(ZFF_X2_fast[12:12]),.I5(ZFF_X2_fast[5:5]),.O(un8_0_8_axb_10));
defparam desc414.INIT=64'h96C33C96693CC369;
  LUT6 un10_axb_10_cZ(.I0(ZFF_Y2[10:10]),.I1(ZFF_Y2[9:9]),.I2(un10_19),.I3(un10_8[15:15]),.I4(un10_8[16:16]),.I5(un10_6[16:16]),.O(un10_axb_10));
defparam un10_axb_10_cZ.INIT=64'hA665599A599AA665;
  LUT5 un10_29_cZ(.I0(ZFF_Y2[10:10]),.I1(ZFF_Y2[9:9]),.I2(un10_19),.I3(un10_8[15:15]),.I4(un10_8[16:16]),.O(un10_29));
defparam un10_29_cZ.INIT=32'hF7755110;
  LUT6 un10_8_axb_16_cZ(.I0(ZFF_Y2_6_rep1),.I1(ZFF_Y2_7_rep1),.I2(ZFF_Y2_8_rep1),.I3(ZFF_Y2[5:5]),.I4(ZFF_Y2[10:10]),.I5(ZFF_Y2[11:11]),.O(un10_8_axb_16));
defparam un10_8_axb_16_cZ.INIT=64'h965AA59669A55A69;
  LUT6 desc415(.I0(ZFF_Y2_fast[7:7]),.I1(ZFF_Y2_fast[6:6]),.I2(ZFF_Y2[12:12]),.I3(ZFF_Y2[10:10]),.I4(ZFF_Y2[11:11]),.I5(ZFF_Y2[13:13]),.O(un10_6_axb_16));
defparam desc415.INIT=64'h95A96A566A5695A9;
  LUT6 desc416(.I0(ZFF_X2_fast[2:2]),.I1(ZFF_X2_fast[10:10]),.I2(ZFF_X2_fast[3:3]),.I3(ZFF_X2_fast[13:13]),.I4(ZFF_X2_fast[11:11]),.I5(ZFF_X2_fast[12:12]),.O(un8_0_8_axb_8));
defparam desc416.INIT=64'hD22D2DD24BB4B44B;
  LUT6 Y_out_double_2_6_0_axb_2_cZ(.I0(pgZFF_X1[1:1]),.I1(pgZFF_X1[2:2]),.I2(pgZFF_Y1[1:1]),.I3(pgZFF_Y1[2:2]),.I4(pgZFF_Y2[1:1]),.I5(pgZFF_Y2[2:2]),.O(Y_out_double_2_6_0_axb_2));
defparam Y_out_double_2_6_0_axb_2_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_15_cZ(.I0(pgZFF_X1[14:14]),.I1(pgZFF_X1[15:15]),.I2(pgZFF_Y1[14:14]),.I3(pgZFF_Y1[15:15]),.I4(pgZFF_Y2[14:14]),.I5(pgZFF_Y2[15:15]),.O(Y_out_double_2_6_0_axb_15));
defparam Y_out_double_2_6_0_axb_15_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_14_cZ(.I0(pgZFF_X1[13:13]),.I1(pgZFF_X1[14:14]),.I2(pgZFF_Y1[13:13]),.I3(pgZFF_Y1[14:14]),.I4(pgZFF_Y2[13:13]),.I5(pgZFF_Y2[14:14]),.O(Y_out_double_2_6_0_axb_14));
defparam Y_out_double_2_6_0_axb_14_cZ.INIT=64'hC639639C39C69C63;
  LUT6 un9_11_s_7_RNI5PQR1(.I0(ZFF_Y1_17_rep1),.I1(un9_11[23:23]),.I2(ZFF_Y1_15_rep1),.I3(un9_11[22:22]),.I4(un9_10[8:8]),.I5(un9_11[28:28]),.O(un9_6_0_axb_28));
defparam un9_11_s_7_RNI5PQR1.INIT=64'h36936339C96C9CC6;
  LUT6 Y_out_double_2_6_0_axb_13_cZ(.I0(pgZFF_X1[12:12]),.I1(pgZFF_X1[13:13]),.I2(pgZFF_Y1[12:12]),.I3(pgZFF_Y1[13:13]),.I4(pgZFF_Y2[12:12]),.I5(pgZFF_Y2[13:13]),.O(Y_out_double_2_6_0_axb_13));
defparam Y_out_double_2_6_0_axb_13_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_12_cZ(.I0(pgZFF_X1[11:11]),.I1(pgZFF_X1[12:12]),.I2(pgZFF_Y1[11:11]),.I3(pgZFF_Y1[12:12]),.I4(pgZFF_Y2[11:11]),.I5(pgZFF_Y2[12:12]),.O(Y_out_double_2_6_0_axb_12));
defparam Y_out_double_2_6_0_axb_12_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_11_cZ(.I0(pgZFF_X1[10:10]),.I1(pgZFF_X1[11:11]),.I2(pgZFF_Y1[10:10]),.I3(pgZFF_Y1[11:11]),.I4(pgZFF_Y2[10:10]),.I5(pgZFF_Y2[11:11]),.O(Y_out_double_2_6_0_axb_11));
defparam Y_out_double_2_6_0_axb_11_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_9_cZ(.I0(pgZFF_X1[8:8]),.I1(pgZFF_X1[9:9]),.I2(pgZFF_Y1[8:8]),.I3(pgZFF_Y1[9:9]),.I4(pgZFF_Y2[8:8]),.I5(pgZFF_Y2[9:9]),.O(Y_out_double_2_6_0_axb_9));
defparam Y_out_double_2_6_0_axb_9_cZ.INIT=64'hC639639C39C69C63;
  LUT5 un8_0_8_axb_11_cZ(.I0(ZFF_X2_fast[15:15]),.I1(ZFF_X2_6_rep1),.I2(ZFF_X2_fast[1:1]),.I3(ZFF_X2_fast[0:0]),.I4(ZFF_X2_fast[5:5]),.O(un8_0_8_axb_11));
defparam un8_0_8_axb_11_cZ.INIT=32'h963CC396;
  LUT6 Y_out_double_2_6_0_axb_7_cZ(.I0(pgZFF_X1[6:6]),.I1(pgZFF_X1[7:7]),.I2(pgZFF_Y1[6:6]),.I3(pgZFF_Y1[7:7]),.I4(pgZFF_Y2[6:6]),.I5(pgZFF_Y2[7:7]),.O(Y_out_double_2_6_0_axb_7));
defparam Y_out_double_2_6_0_axb_7_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_6_cZ(.I0(pgZFF_X1[5:5]),.I1(pgZFF_X1[6:6]),.I2(pgZFF_Y1[5:5]),.I3(pgZFF_Y1[6:6]),.I4(pgZFF_Y2[5:5]),.I5(pgZFF_Y2[6:6]),.O(Y_out_double_2_6_0_axb_6));
defparam Y_out_double_2_6_0_axb_6_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_5_cZ(.I0(pgZFF_X1[4:4]),.I1(pgZFF_X1[5:5]),.I2(pgZFF_Y1[4:4]),.I3(pgZFF_Y1[5:5]),.I4(pgZFF_Y2[4:4]),.I5(pgZFF_Y2[5:5]),.O(Y_out_double_2_6_0_axb_5));
defparam Y_out_double_2_6_0_axb_5_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_3_cZ(.I0(pgZFF_X1[2:2]),.I1(pgZFF_X1[3:3]),.I2(pgZFF_Y1[2:2]),.I3(pgZFF_Y1[3:3]),.I4(pgZFF_Y2[2:2]),.I5(pgZFF_Y2[3:3]),.O(Y_out_double_2_6_0_axb_3));
defparam Y_out_double_2_6_0_axb_3_cZ.INIT=64'hC639639C39C69C63;
  LUT5 un9_8_axb_14_cZ(.I0(ZFF_Y1_fast[17:17]),.I1(ZFF_Y1_fast[7:7]),.I2(un9_8_6_rep1),.I3(ZFF_Y1_fast[8:8]),.I4(un9_10_8_rep1),.O(un9_8_axb_14));
defparam un9_8_axb_14_cZ.INIT=32'h78871EE1;
  LUT6 un9_axb_8_cZ(.I0(ZFF_Y1[7:7]),.I1(ZFF_Y1[5:5]),.I2(un9_8[9:9]),.I3(un9_8[10:10]),.I4(un9_6[10:10]),.I5(un9_6[9:9]),.O(un9_axb_8));
defparam un9_axb_8_cZ.INIT=64'h39C6C6399C63639C;
  LUT6 un7_0_0_axb_17_cZ(.I0(ZFF_X1[13:13]),.I1(un7_0_10_i_i[17:17]),.I2(un7_0_6[17:17]),.I3(un7_0_6[16:16]),.I4(un7_0_8[17:17]),.I5(un7_0_8[16:16]),.O(un7_0_0_axb_17));
defparam un7_0_0_axb_17_cZ.INIT=64'h3C69C39669C3963C;
  LUT6 un10_axb_18_cZ(.I0(ZFF_Y2[16:16]),.I1(ZFF_Y2[15:15]),.I2(un10_8[23:23]),.I3(un10_8[24:24]),.I4(un10_6[23:23]),.I5(un10_6[24:24]),.O(un10_axb_18));
defparam un10_axb_18_cZ.INIT=64'hA659659A59A69A65;
  LUT6 un10_8_axb_21_cZ(.I0(ZFF_Y2[12:12]),.I1(ZFF_Y2[10:10]),.I2(ZFF_Y2[11:11]),.I3(ZFF_Y2[13:13]),.I4(ZFF_Y2[16:16]),.I5(ZFF_Y2[15:15]),.O(un10_8_axb_21));
defparam un10_8_axb_21_cZ.INIT=64'h87787887E11E1EE1;
  LUT6 un10_axb_16_cZ(.I0(ZFF_Y2[16:16]),.I1(ZFF_Y2[15:15]),.I2(un10_8[21:21]),.I3(un10_8[22:22]),.I4(un10_6[21:21]),.I5(un10_6[22:22]),.O(un10_axb_16));
defparam un10_axb_16_cZ.INIT=64'hA659659A59A69A65;
  LUT6 desc417(.I0(ZFF_Y2_fast[8:8]),.I1(ZFF_Y2[5:5]),.I2(ZFF_Y2[0:0]),.I3(ZFF_Y2[2:2]),.I4(ZFF_Y2[1:1]),.I5(ZFF_Y2[13:13]),.O(un10_6_axb_5));
defparam desc417.INIT=64'h5AA596699669A55A;
  LUT6 desc418(.I0(ZFF_Y2_fast[7:7]),.I1(ZFF_Y2_fast[6:6]),.I2(ZFF_Y2_8_rep1),.I3(ZFF_Y2[5:5]),.I4(ZFF_Y2[2:2]),.I5(ZFF_Y2[1:1]),.O(un10_6_axb_11));
defparam desc418.INIT=64'h96C3693C3C96C369;
  LUT6 ZFF_X2_6_rep1_RNIRKED1(.I0(ZFF_X2_6_rep1),.I1(ZFF_X2_2_rep1),.I2(ZFF_X2_fast[1:1]),.I3(ZFF_X2_fast[0:0]),.I4(ZFF_X2_fast[12:12]),.I5(ZFF_X2[11:11]),.O(un8_0_6_axb_7));
defparam ZFF_X2_6_rep1_RNIRKED1.INIT=64'h936C6C93C93636C9;
  LUT5 desc419(.I0(ZFF_X1[3:3]),.I1(ZFF_X1_fast[16:16]),.I2(ZFF_X1[4:4]),.I3(ZFF_X1[6:6]),.I4(ZFF_X1[7:7]),.O(un7_0_10_axb_14));
defparam desc419.INIT=32'hB4D24B2D;
  LUT5 desc420(.I0(ZFF_X1_fast[12:12]),.I1(ZFF_X1_fast[13:13]),.I2(ZFF_X1_fast[3:3]),.I3(ZFF_X1_fast[2:2]),.I4(ZFF_X1_fast[4:4]),.O(un7_0_6_axb_10));
defparam desc420.INIT=32'hC96C3693;
  LUT6 ZFF_Y2_14_rep1_RNIUGK11(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2[10:10]),.I2(ZFF_Y2[13:13]),.I3(ZFF_Y2[16:16]),.I4(ZFF_Y2[15:15]),.I5(ZFF_Y2[9:9]),.O(un10_6_axb_19));
defparam ZFF_Y2_14_rep1_RNIUGK11.INIT=64'h9966699669966699;
  LUT6 un10_8_axb_19_cZ(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2_8_rep1),.I2(ZFF_Y2[10:10]),.I3(ZFF_Y2[11:11]),.I4(ZFF_Y2[13:13]),.I5(ZFF_Y2[9:9]),.O(un10_8_axb_19));
defparam un10_8_axb_19_cZ.INIT=64'h956AA9566A9556A9;
  LUT6 un10_axb_14_cZ(.I0(ZFF_Y2[14:14]),.I1(ZFF_Y2[13:13]),.I2(un10_8[19:19]),.I3(un10_8[20:20]),.I4(un10_6[19:19]),.I5(un10_6[20:20]),.O(un10_axb_14));
defparam un10_axb_14_cZ.INIT=64'hA659659A59A69A65;
  LUT6 ZFF_X0_11_rep1_RNIFACJ1(.I0(ZFF_X0_11_rep1),.I1(ZFF_X0_6_rep1),.I2(ZFF_X0_2_rep1),.I3(ZFF_X0_12_rep1),.I4(ZFF_X0_fast[0:0]),.I5(ZFF_X0_1_rep1),.O(un6_0_6_axb_7));
defparam ZFF_X0_11_rep1_RNIFACJ1.INIT=64'hD22D2DD24BB4B44B;
  LUT5 Y_out_double_2_6_0_axb_17_cZ(.I0(pgZFF_Y1[17:17]),.I1(pgZFF_Y2[17:17]),.I2(pgZFF_X1[17:17]),.I3(pgZFF_Y1[16:16]),.I4(pgZFF_Y2[16:16]),.O(Y_out_double_2_6_0_axb_17));
defparam Y_out_double_2_6_0_axb_17_cZ.INIT=32'h96666669;
  LUT6 Y_out_double_2_6_0_axb_16_cZ(.I0(pgZFF_X1[17:17]),.I1(pgZFF_Y1[16:16]),.I2(pgZFF_Y2[16:16]),.I3(pgZFF_X1[15:15]),.I4(pgZFF_Y1[15:15]),.I5(pgZFF_Y2[15:15]),.O(Y_out_double_2_6_0_axb_16));
defparam Y_out_double_2_6_0_axb_16_cZ.INIT=64'h9696699669966969;
  LUT6 desc421(.I0(ZFF_X0_fast[14:14]),.I1(ZFF_X0_fast[15:15]),.I2(ZFF_X0_fast[12:12]),.I3(ZFF_X0_fast[4:4]),.I4(ZFF_X0_fast[0:0]),.I5(ZFF_X0_fast[5:5]),.O(un6_0_8_axb_10));
defparam desc421.INIT=64'h93C96C366C3693C9;
  LUT6 desc422(.I0(ZFF_X0_fast[2:2]),.I1(ZFF_X0_fast[10:10]),.I2(ZFF_X0_fast[12:12]),.I3(ZFF_X0_fast[11:11]),.I4(ZFF_X0_fast[3:3]),.I5(ZFF_X0_fast[13:13]),.O(un6_0_8_axb_8));
defparam desc422.INIT=64'hD42B2BD42BD4D42B;
  LUT6 Y_out_double_2_6_0_axb_10_cZ(.I0(pgZFF_X1[9:9]),.I1(pgZFF_X1[10:10]),.I2(pgZFF_Y1[9:9]),.I3(pgZFF_Y1[10:10]),.I4(pgZFF_Y2[9:9]),.I5(pgZFF_Y2[10:10]),.O(Y_out_double_2_6_0_axb_10));
defparam Y_out_double_2_6_0_axb_10_cZ.INIT=64'hC639639C39C69C63;
  LUT6 Y_out_double_2_6_0_axb_8_cZ(.I0(pgZFF_X1[7:7]),.I1(pgZFF_X1[8:8]),.I2(pgZFF_Y1[7:7]),.I3(pgZFF_Y1[8:8]),.I4(pgZFF_Y2[7:7]),.I5(pgZFF_Y2[8:8]),.O(Y_out_double_2_6_0_axb_8));
defparam Y_out_double_2_6_0_axb_8_cZ.INIT=64'hC639639C39C69C63;
  LUT6 desc423(.I0(ZFF_X2_fast[14:14]),.I1(ZFF_X2_fast[3:3]),.I2(ZFF_X2_fast[13:13]),.I3(ZFF_X2_fast[11:11]),.I4(ZFF_X2_fast[4:4]),.I5(ZFF_X2_fast[12:12]),.O(un8_0_8_axb_9));
defparam desc423.INIT=64'hA665599A599AA665;
  LUT6 desc424(.I0(ZFF_X2_fast[2:2]),.I1(ZFF_X2_fast[10:10]),.I2(ZFF_X2_fast[1:1]),.I3(ZFF_X2_fast[11:11]),.I4(ZFF_X2_fast[12:12]),.I5(ZFF_X2_fast[9:9]),.O(un8_0_8_axb_7));
defparam desc424.INIT=64'h9969669669669699;
  LUT6 Y_out_double_2_6_0_axb_4_cZ(.I0(pgZFF_X1[3:3]),.I1(pgZFF_X1[4:4]),.I2(pgZFF_Y1[3:3]),.I3(pgZFF_Y1[4:4]),.I4(pgZFF_Y2[3:3]),.I5(pgZFF_Y2[4:4]),.O(Y_out_double_2_6_0_axb_4));
defparam Y_out_double_2_6_0_axb_4_cZ.INIT=64'hC639639C39C69C63;
  LUT6 un10_8_axb_17_cZ(.I0(ZFF_Y2_6_rep1),.I1(ZFF_Y2_7_rep1),.I2(ZFF_Y2_8_rep1),.I3(ZFF_Y2[12:12]),.I4(ZFF_Y2[11:11]),.I5(ZFF_Y2[9:9]),.O(un10_8_axb_17));
defparam un10_8_axb_17_cZ.INIT=64'h936CC9366C9336C9;
  LUT6 ZFF_Y2_7_rep1_RNI7K501(.I0(ZFF_Y2_7_rep1),.I1(ZFF_Y2_14_rep1),.I2(ZFF_Y2_8_rep1),.I3(ZFF_Y2[12:12]),.I4(ZFF_Y2[11:11]),.I5(ZFF_Y2[13:13]),.O(un10_6_axb_17));
defparam ZFF_Y2_7_rep1_RNI7K501.INIT=64'h9669C33C3CC39669;
  LUT6 un10_axb_12_cZ(.I0(ZFF_Y2[12:12]),.I1(ZFF_Y2[11:11]),.I2(un10_8[17:17]),.I3(un10_29),.I4(un10_8[18:18]),.I5(un10_6[18:18]),.O(un10_axb_12));
defparam un10_axb_12_cZ.INIT=64'hA665599A599AA665;
  LUT6 desc425(.I0(un9_11_fast[26:26]),.I1(un9_8_fast[7:7]),.I2(un9_8_fast[6:6]),.I3(ZFF_Y1_fast[5:5]),.I4(un9_11_fast[25:25]),.I5(ZFF_Y1_fast[6:6]),.O(un9_8_axb_8));
defparam desc425.INIT=64'h9699669669669969;
  LUT5 un9_8_axb_18_cZ(.I0(un9_11_fast[24:24]),.I1(ZFF_Y1_17_rep1),.I2(un9_11_fast[23:23]),.I3(ZFF_Y1_5_rep1),.I4(ZFF_Y1_4_rep1),.O(un9_8_axb_18));
defparam un9_8_axb_18_cZ.INIT=32'h6A9556A9;
  LUT6 un9_11_axb_6_RNILUBQ(.I0(ZFF_Y1_17_rep1),.I1(ZFF_Y1_9_rep1),.I2(un9_11_26_rep1),.I3(ZFF_Y1_16_rep1),.I4(un9_11[22:22]),.I5(un9_11[27:27]),.O(un9_6_0_axb_27));
defparam un9_11_axb_6_RNILUBQ.INIT=64'h566AA995A995566A;
  LUT6 un10_axb_15_cZ(.I0(ZFF_Y2[14:14]),.I1(ZFF_Y2[15:15]),.I2(un10_8[20:20]),.I3(un10_8[21:21]),.I4(un10_6[20:20]),.I5(un10_6[21:21]),.O(un10_axb_15));
defparam un10_axb_15_cZ.INIT=64'hC639639C39C69C63;
  LUT6 un10_8_axb_20_cZ(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2[12:12]),.I2(ZFF_Y2[10:10]),.I3(ZFF_Y2[11:11]),.I4(ZFF_Y2[15:15]),.I5(ZFF_Y2[9:9]),.O(un10_8_axb_20));
defparam un10_8_axb_20_cZ.INIT=64'hC3693C96693C96C3;
  LUT6 un9_axb_36_cZ(.I0(un9_8[37:37]),.I1(un9_10[37:37]),.I2(un9_10[38:38]),.I3(un9_8[38:38]),.I4(un9_6[37:37]),.I5(un9_6[38:38]),.O(un9_axb_36));
defparam un9_axb_36_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 un10_8_axb_15_cZ(.I0(ZFF_Y2_6_rep1),.I1(ZFF_Y2_7_rep1),.I2(ZFF_Y2[4:4]),.I3(ZFF_Y2[5:5]),.I4(ZFF_Y2[10:10]),.I5(ZFF_Y2[9:9]),.O(un10_8_axb_15));
defparam un10_8_axb_15_cZ.INIT=64'h936C6C93C93636C9;
  LUT6 desc426(.I0(ZFF_Y2_fast[6:6]),.I1(ZFF_Y2[5:5]),.I2(ZFF_Y2[12:12]),.I3(ZFF_Y2[10:10]),.I4(ZFF_Y2[11:11]),.I5(ZFF_Y2[9:9]),.O(un10_6_axb_15));
defparam desc426.INIT=64'h96695AA5A55A9669;
  LUT6 desc427(.I0(ZFF_Y2_fast[6:6]),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[5:5]),.I3(ZFF_Y2[0:0]),.I4(ZFF_Y2[3:3]),.I5(ZFF_Y2[9:9]),.O(un10_6_axb_9));
defparam desc427.INIT=64'h6699966996699966;
  LUT6 ZFF_Y2_8_rep1_RNIBDPL1(.I0(ZFF_Y2_8_rep1),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[5:5]),.I3(ZFF_Y2[10:10]),.I4(ZFF_Y2[11:11]),.I5(ZFF_Y2[9:9]),.O(un10_6_axb_14));
defparam ZFF_Y2_8_rep1_RNIBDPL1.INIT=64'hD24B2DB42DB4D24B;
  LUT6 un10_8_axb_14_cZ(.I0(ZFF_Y2_6_rep1),.I1(ZFF_Y2_8_rep1),.I2(ZFF_Y2[4:4]),.I3(ZFF_Y2[5:5]),.I4(ZFF_Y2[3:3]),.I5(ZFF_Y2[9:9]),.O(un10_8_axb_14));
defparam un10_8_axb_14_cZ.INIT=64'hA569695A5A9696A5;
  LUT6 desc428(.I0(ZFF_Y2_fast[8:8]),.I1(ZFF_Y2[0:0]),.I2(ZFF_Y2[3:3]),.I3(ZFF_Y2[2:2]),.I4(ZFF_Y2[1:1]),.I5(ZFF_Y2[15:15]),.O(un10_6_axb_6));
defparam desc428.INIT=64'h781E87E187E1781E;
  LUT6 un10_8_axb_13_cZ(.I0(ZFF_Y2_7_rep1),.I1(ZFF_Y2_8_rep1),.I2(ZFF_Y2[4:4]),.I3(ZFF_Y2[5:5]),.I4(ZFF_Y2[3:3]),.I5(ZFF_Y2[2:2]),.O(un10_8_axb_13));
defparam un10_8_axb_13_cZ.INIT=64'hC63939C6639C9C63;
  LUT6 desc429(.I0(ZFF_Y2_fast[7:7]),.I1(ZFF_Y2_8_rep1),.I2(ZFF_Y2[4:4]),.I3(ZFF_Y2[3:3]),.I4(ZFF_Y2[10:10]),.I5(ZFF_Y2[9:9]),.O(un10_6_axb_13));
defparam desc429.INIT=64'hC3693C96693C96C3;
  LUT6 un10_8_axb_12_cZ(.I0(ZFF_Y2_6_rep1),.I1(ZFF_Y2_7_rep1),.I2(ZFF_Y2[4:4]),.I3(ZFF_Y2[3:3]),.I4(ZFF_Y2[2:2]),.I5(ZFF_Y2[1:1]),.O(un10_8_axb_12));
defparam un10_8_axb_12_cZ.INIT=64'hC3693C96693C96C3;
  LUT6 desc430(.I0(ZFF_Y2_fast[7:7]),.I1(ZFF_Y2_fast[6:6]),.I2(ZFF_Y2_8_rep1),.I3(ZFF_Y2[3:3]),.I4(ZFF_Y2[2:2]),.I5(ZFF_Y2[9:9]),.O(un10_6_axb_12));
defparam desc430.INIT=64'hA659659A59A69A65;
  LUT6 desc431(.I0(ZFF_X1_fast[15:15]),.I1(ZFF_X1_fast[9:9]),.I2(ZFF_X1_fast[5:5]),.I3(ZFF_X1_fast[8:8]),.I4(ZFF_X1_fast[4:4]),.I5(ZFF_X1_fast[14:14]),.O(un7_0_6_axb_12));
defparam desc431.INIT=64'h9669696996969669;
  LUT6 un10_axb_19_cZ(.I0(ZFF_Y2[16:16]),.I1(ZFF_Y2[17:17]),.I2(un10_8[24:24]),.I3(un10_8[25:25]),.I4(un10_6[24:24]),.I5(un10_6[25:25]),.O(un10_axb_19));
defparam un10_axb_19_cZ.INIT=64'hC639639C39C69C63;
  LUT6 un10_axb_17_cZ(.I0(ZFF_Y2[16:16]),.I1(ZFF_Y2[15:15]),.I2(un10_8[22:22]),.I3(un10_8[23:23]),.I4(un10_6[22:22]),.I5(un10_6[23:23]),.O(un10_axb_17));
defparam un10_axb_17_cZ.INIT=64'hC639639C39C69C63;
  LUT6 un10_8_axb_22_cZ(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2[12:12]),.I2(ZFF_Y2[11:11]),.I3(ZFF_Y2[13:13]),.I4(ZFF_Y2[16:16]),.I5(ZFF_Y2[17:17]),.O(un10_8_axb_22));
defparam un10_8_axb_22_cZ.INIT=64'h9666999669996669;
  LUT6 un10_8_axb_18_cZ(.I0(ZFF_Y2_7_rep1),.I1(ZFF_Y2_8_rep1),.I2(ZFF_Y2[12:12]),.I3(ZFF_Y2[10:10]),.I4(ZFF_Y2[13:13]),.I5(ZFF_Y2[9:9]),.O(un10_8_axb_18));
defparam un10_8_axb_18_cZ.INIT=64'h9C63639C39C6C639;
  LUT6 ZFF_Y2_14_rep1_RNIF2RA1(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2_8_rep1),.I2(ZFF_Y2[12:12]),.I3(ZFF_Y2[13:13]),.I4(ZFF_Y2[15:15]),.I5(ZFF_Y2[9:9]),.O(un10_6_axb_18));
defparam ZFF_Y2_14_rep1_RNIF2RA1.INIT=64'h8E71718E718E8E71;
  LUT6 un10_axb_13_cZ(.I0(ZFF_Y2[12:12]),.I1(ZFF_Y2[13:13]),.I2(un10_8[18:18]),.I3(un10_8[19:19]),.I4(un10_6[18:18]),.I5(un10_6[19:19]),.O(un10_axb_13));
defparam un10_axb_13_cZ.INIT=64'hC639639C39C69C63;
  LUT5 desc432(.I0(ZFF_X1_fast[13:13]),.I1(ZFF_X1_fast[3:3]),.I2(ZFF_X1_fast[8:8]),.I3(ZFF_X1_fast[4:4]),.I4(ZFF_X1_fast[14:14]),.O(un7_0_6_axb_11));
defparam desc432.INIT=32'hD2B42D4B;
  LUT6 desc433(.I0(ZFF_X1_fast[15:15]),.I1(ZFF_X1_fast[9:9]),.I2(ZFF_X1_fast[10:10]),.I3(ZFF_X1_fast[5:5]),.I4(ZFF_X1_fast[6:6]),.I5(ZFF_X1_fast[16:16]),.O(un7_0_6_axb_13));
defparam desc433.INIT=64'hD24B2DB42DB4D24B;
  LUT5 un10_axb_23_cZ(.I0(ZFF_Y2[17:17]),.I1(un10_8[28:28]),.I2(un10_8[29:29]),.I3(un10_6[28:28]),.I4(un10_6[29:29]),.O(un10_axb_23));
defparam un10_axb_23_cZ.INIT=32'h2DB4D24B;
  LUT4 un9_o5_36_cZ(.I0(ZFF_Y1[16:16]),.I1(un9_8_cry_29),.I2(un9_10[38:38]),.I3(un9_6[38:38]),.O(un9_o5_36));
defparam un9_o5_36_cZ.INIT=16'hF990;
  LUT6 desc434(.I0(ZFF_Y1_fast[16:16]),.I1(un9_11_fast[26:26]),.I2(ZFF_Y1_fast[4:4]),.I3(un9_11_fast[22:22]),.I4(ZFF_Y1_fast[5:5]),.I5(ZFF_Y1_fast[9:9]),.O(un9_8_axb_11));
defparam desc434.INIT=64'h6C3693C993C96C36;
  LUT5 un9_axb_10_cZ(.I0(un9_8[7:7]),.I1(un9_10[8:8]),.I2(un9_8[12:12]),.I3(un9_6[12:12]),.I4(un9_o5_9),.O(un9_axb_10));
defparam un9_axb_10_cZ.INIT=32'h96696996;
  LUT5 ZFF_X1_1_rep1_RNIQ69J1(.I0(ZFF_X1_1_rep1),.I1(ZFF_X1_0_rep1),.I2(ZFF_X1_7_rep1),.I3(ZFF_X1_8_rep1),.I4(ZFF_X1_fast[16:16]),.O(un7_0_6_axb_15));
defparam ZFF_X1_1_rep1_RNIQ69J1.INIT=32'h9A65A659;
  LUT6 ZFF_Y1_8_rep1_RNI1S771(.I0(ZFF_Y1_8_rep1),.I1(ZFF_Y1_9_rep1),.I2(ZFF_Y1_6_rep1),.I3(ZFF_Y1_3_rep1),.I4(ZFF_Y1_5_rep1),.I5(un9_8[7:7]),.O(un9_10_axb_16));
defparam ZFF_Y1_8_rep1_RNI1S771.INIT=64'h3CC369966996C33C;
  LUT6 ZFF_Y1_9_rep1_RNIK1602(.I0(ZFF_Y1_9_rep1),.I1(ZFF_Y1[4:4]),.I2(ZFF_Y1[6:6]),.I3(ZFF_Y1_7_rep1),.I4(un9_11[22:22]),.I5(ZFF_Y1[3:3]),.O(un9_10_axb_17));
defparam ZFF_Y1_9_rep1_RNIK1602.INIT=64'h36C9C9366C93936C;
  LUT6 ZFF_X2_14_rep1_RNILLJ61(.I0(ZFF_X2_14_rep1),.I1(ZFF_X2[10:10]),.I2(ZFF_X2[9:9]),.I3(ZFF_X2[8:8]),.I4(ZFF_X2[11:11]),.I5(ZFF_X2_fast[16:16]),.O(un8_0_6_axb_16));
defparam ZFF_X2_14_rep1_RNILLJ61.INIT=64'h69A5965A5A69A596;
  LUT6 un10_axb_5_cZ(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[5:5]),.I3(ZFF_Y2[3:3]),.I4(ZFF_Y2[1:1]),.I5(un10_6[11:11]),.O(un10_axb_5));
defparam un10_axb_5_cZ.INIT=64'hF0F0F0D20F0F0F2D;
  LUT6 un6_0_0_axb_17_cZ(.I0(un6_0_8[16:16]),.I1(un6_0_8[17:17]),.I2(un6_0_9[16:16]),.I3(un6_0_9[17:17]),.I4(un6_0_6[16:16]),.I5(un6_0_6[17:17]),.O(un6_0_0_axb_17));
defparam un6_0_0_axb_17_cZ.INIT=64'h36C96C93C936936C;
  LUT6 desc435(.I0(un9_11_fast[26:26]),.I1(un9_11_22_rep1),.I2(ZFF_Y1_6_rep1),.I3(un9_11_23_rep1),.I4(ZFF_Y1_5_rep1),.I5(ZFF_Y1_15_rep1),.O(un9_6_0_axb_23));
defparam desc435.INIT=64'h1EE17887E11E8778;
  LUT5 desc436(.I0(ZFF_X2_fast[6:6]),.I1(ZFF_X2_fast[8:8]),.I2(ZFF_X2_fast[4:4]),.I3(ZFF_X2_fast[7:7]),.I4(ZFF_X2_fast[5:5]),.O(un8_0_8_axb_3));
defparam desc436.INIT=32'h66699666;
  LUT6 desc437(.I0(ZFF_X1_fast[12:12]),.I1(ZFF_X1_fast[13:13]),.I2(ZFF_X1_4_rep1),.I3(ZFF_X1_fast[5:5]),.I4(ZFF_X1_6_rep1),.I5(ZFF_X1_7_rep1),.O(un7_0_8_axb_10));
defparam desc437.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_15_cZ(.I0(ZFF_X0[7:7]),.I1(ZFF_X0[8:8]),.I2(un6_0_8[14:14]),.I3(un6_0_8[15:15]),.I4(un6_0_6[14:14]),.I5(un6_0_6[15:15]),.O(un6_0_0_axb_15));
defparam un6_0_0_axb_15_cZ.INIT=64'h9669669969969966;
  LUT3 un10_o5_12_cZ(.I0(ZFF_Y2[12:12]),.I1(un10_8[18:18]),.I2(un10_6[18:18]),.O(un10_o5_12));
defparam un10_o5_12_cZ.INIT=8'hD4;
  LUT6 ZFF_X2_15_rep1_RNIKV8G1(.I0(ZFF_X2_15_rep1),.I1(ZFF_X2[3:3]),.I2(ZFF_X2[4:4]),.I3(ZFF_X2[6:6]),.I4(ZFF_X2[5:5]),.I5(ZFF_X2_fast[16:16]),.O(un8_0_6_axb_11));
defparam ZFF_X2_15_rep1_RNIKV8G1.INIT=64'hD22D4BB42DD2B44B;
  LUT5 desc438(.I0(ZFF_X2_fast[6:6]),.I1(ZFF_X2_fast[8:8]),.I2(ZFF_X2_fast[7:7]),.I3(ZFF_X2_fast[9:9]),.I4(ZFF_X2_fast[5:5]),.O(un8_0_8_axb_4));
defparam desc438.INIT=32'h4BB42DD2;
  LUT3 un10_8_o5_17_cZ(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[12:12]),.I2(ZFF_Y2[9:9]),.O(un10_8_o5_17));
defparam un10_8_o5_17_cZ.INIT=8'hB2;
  LUT3 un10_8_o5_18_cZ(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[10:10]),.I2(ZFF_Y2[13:13]),.O(un10_8_o5_18));
defparam un10_8_o5_18_cZ.INIT=8'h8E;
  LUT6 desc439(.I0(ZFF_X1_fast[13:13]),.I1(ZFF_X1_fast[5:5]),.I2(ZFF_X1_6_rep1),.I3(ZFF_X1_7_rep1),.I4(ZFF_X1_fast[14:14]),.I5(ZFF_X1_8_rep1),.O(un7_0_8_axb_11));
defparam desc439.INIT=64'h1E78E187E1871E78;
  LUT5 desc440(.I0(ZFF_X1[3:3]),.I1(ZFF_X1[2:2]),.I2(ZFF_X1[5:5]),.I3(ZFF_X1_fast[16:16]),.I4(ZFF_X1[6:6]),.O(un7_0_10_axb_13));
defparam desc440.INIT=32'h59A6A659;
  LUT5 desc441(.I0(ZFF_X2_fast[10:10]),.I1(ZFF_X2_fast[1:1]),.I2(ZFF_X2_fast[11:11]),.I3(ZFF_X2_fast[0:0]),.I4(ZFF_X2_fast[9:9]),.O(un8_0_8_axb_6));
defparam desc441.INIT=32'h96C3693C;
  LUT6 ZFF_X0_14_rep1_RNI4VP72(.I0(ZFF_X0_14_rep1),.I1(ZFF_X0_15_rep1),.I2(ZFF_X0[10:10]),.I3(ZFF_X0[9:9]),.I4(ZFF_X0[12:12]),.I5(ZFF_X0[11:11]),.O(un6_0_6_axb_17));
defparam ZFF_X0_14_rep1_RNI4VP72.INIT=64'h3C69C39669C3963C;
  LUT5 ZFF_X0_10_rep1_RNICIH81(.I0(ZFF_X0_10_rep1),.I1(ZFF_X0_14_rep1),.I2(ZFF_X0_15_rep1),.I3(ZFF_X0_fast[16:16]),.I4(ZFF_X0[9:9]),.O(un6_0_8_axb_20));
defparam ZFF_X0_10_rep1_RNICIH81.INIT=32'hA59669A5;
  LUT6 ZFF_X1_4_rep1_RNISEAL1(.I0(ZFF_X1_4_rep1),.I1(ZFF_X1_12_rep1),.I2(ZFF_X1_3_rep1),.I3(ZFF_X1_11_rep1),.I4(ZFF_X1_13_rep1),.I5(ZFF_X1_fast[14:14]),.O(un7_0_8_axb_17));
defparam ZFF_X1_4_rep1_RNISEAL1.INIT=64'h6669699999969666;
  LUT6 ZFF_Y1_11_rep1_RNI1JK02(.I0(un9_11_23_rep1),.I1(ZFF_Y1[5:5]),.I2(ZFF_Y1[4:4]),.I3(ZFF_Y1[8:8]),.I4(ZFF_Y1_7_rep1),.I5(un9_11[22:22]),.O(un9_10_axb_18));
defparam ZFF_Y1_11_rep1_RNI1JK02.INIT=64'h6699699669969966;
  LUT6 un7_0_0_axb_15_cZ(.I0(ZFF_X1[12:12]),.I1(ZFF_X1[11:11]),.I2(un7_0_6[14:14]),.I3(un7_0_6[15:15]),.I4(un7_0_8[14:14]),.I5(un7_0_8[15:15]),.O(un7_0_0_axb_15));
defparam un7_0_0_axb_15_cZ.INIT=64'h56A96A95A956956A;
  LUT6 ZFF_X0_4_rep1_RNIDI4G1(.I0(ZFF_X0_2_rep1),.I1(ZFF_X0_4_rep1),.I2(ZFF_X0_3_rep1),.I3(ZFF_X0_14_rep1),.I4(ZFF_X0_15_rep1),.I5(ZFF_X0[5:5]),.O(un6_0_6_axb_10));
defparam ZFF_X0_4_rep1_RNIDI4G1.INIT=64'h87E1781E781E87E1;
  LUT5 desc442(.I0(ZFF_X0_fast[3:3]),.I1(ZFF_X0_7_rep1),.I2(ZFF_X0_2_rep1),.I3(ZFF_X0_fast[8:8]),.I4(ZFF_X0_fast[16:16]),.O(un6_0_8_axb_13));
defparam desc442.INIT=32'hA65959A6;
  LUT3 un10_o5_14_cZ(.I0(ZFF_Y2[14:14]),.I1(un10_8[20:20]),.I2(un10_6[20:20]),.O(un10_o5_14));
defparam un10_o5_14_cZ.INIT=8'hD4;
  LUT6 un7_0_0_axb_16_cZ(.I0(ZFF_X1[13:13]),.I1(ZFF_X1[12:12]),.I2(un7_0_6[15:15]),.I3(un7_0_6[16:16]),.I4(un7_0_8[15:15]),.I5(un7_0_8[16:16]),.O(un7_0_0_axb_16));
defparam un7_0_0_axb_16_cZ.INIT=64'h56A96A95A956956A;
  LUT3 un8_0_8_o5_10_cZ(.I0(ZFF_X2_fast[15:15]),.I1(ZFF_X2_fast[0:0]),.I2(ZFF_X2_fast[5:5]),.O(un8_0_8_o5_10));
defparam un8_0_8_o5_10_cZ.INIT=8'h8E;
  LUT6 ZFF_X1_4_rep1_RNI2D731(.I0(ZFF_X1_4_rep1),.I1(ZFF_X1_12_rep1),.I2(ZFF_X1_5_rep1),.I3(ZFF_X1_13_rep1),.I4(ZFF_X1_15_rep1),.I5(ZFF_X1_fast[14:14]),.O(un7_0_8_axb_18));
defparam ZFF_X1_4_rep1_RNI2D731.INIT=64'h1EE1E11E78878778;
  LUT6 ZFF_X0_6_rep1_RNIJG1E1(.I0(ZFF_X0_6_rep1),.I1(ZFF_X0_4_rep1),.I2(ZFF_X0_3_rep1),.I3(ZFF_X0_16_rep1),.I4(ZFF_X0_15_rep1),.I5(ZFF_X0[5:5]),.O(un6_0_6_axb_11));
defparam ZFF_X0_6_rep1_RNIJG1E1.INIT=64'h9669996666999669;
  LUT3 un10_8_o5_13_cZ(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[5:5]),.I2(ZFF_Y2[3:3]),.O(un10_8_o5_13));
defparam un10_8_o5_13_cZ.INIT=8'hD4;
  LUT5 desc443(.I0(ZFF_X2[4:4]),.I1(ZFF_X2[6:6]),.I2(ZFF_X2[5:5]),.I3(ZFF_X2[7:7]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_6_axb_12));
defparam desc443.INIT=32'h87781EE1;
  LUT6 desc444(.I0(ZFF_Y2[4:4]),.I1(ZFF_Y2[5:5]),.I2(ZFF_Y2[0:0]),.I3(ZFF_Y2[12:12]),.I4(ZFF_Y2[1:1]),.I5(ZFF_Y2[13:13]),.O(un10_6_axb_4));
defparam desc444.INIT=64'hC663399C399CC663;
  LUT6 ZFF_X0_14_rep1_RNIQUVN1(.I0(ZFF_X0_14_rep1),.I1(ZFF_X0_16_rep1),.I2(ZFF_X0[10:10]),.I3(ZFF_X0[9:9]),.I4(ZFF_X0[8:8]),.I5(ZFF_X0[11:11]),.O(un6_0_6_axb_16));
defparam ZFF_X0_14_rep1_RNIQUVN1.INIT=64'h59A69A65A659659A;
  LUT6 ZFF_X2_2_rep1_RNIIIMJ1(.I0(ZFF_X2_2_rep1),.I1(ZFF_X2_10_rep1),.I2(ZFF_X2_fast[0:0]),.I3(ZFF_X2_fast[4:4]),.I4(ZFF_X2_fast[5:5]),.I5(ZFF_X2[9:9]),.O(un8_0_6_axb_5));
defparam ZFF_X2_2_rep1_RNIIIMJ1.INIT=64'h963C69C3C3963C69;
  LUT5 desc445(.I0(ZFF_X0_fast[7:7]),.I1(ZFF_X0_fast[6:6]),.I2(ZFF_X0_fast[9:9]),.I3(ZFF_X0_fast[8:8]),.I4(ZFF_X0_fast[5:5]),.O(un6_0_8_axb_4));
defparam desc445.INIT=32'h695A5A96;
  LUT5 ZFF_X0_16_rep1_RNI7TU91(.I0(ZFF_X0_16_rep1),.I1(ZFF_X0[7:7]),.I2(ZFF_X0[10:10]),.I3(ZFF_X0[9:9]),.I4(ZFF_X0[8:8]),.O(un6_0_6_axb_15));
defparam ZFF_X0_16_rep1_RNI7TU91.INIT=32'h871E78E1;
  LUT6 un6_0_0_axb_19_cZ(.I0(un6_0_8[18:18]),.I1(un6_0_8[19:19]),.I2(un6_0_9[18:18]),.I3(un6_0_9[19:19]),.I4(un6_0_6[18:18]),.I5(un6_0_6[19:19]),.O(un6_0_0_axb_19));
defparam un6_0_0_axb_19_cZ.INIT=64'h36C96C93C936936C;
  LUT3 un10_8_o5_16_cZ(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[6:6]),.I2(ZFF_Y2[11:11]),.O(un10_8_o5_16));
defparam un10_8_o5_16_cZ.INIT=8'h8E;
  LUT3 un10_8_o5_14_cZ(.I0(ZFF_Y2[6:6]),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[9:9]),.O(un10_8_o5_14));
defparam un10_8_o5_14_cZ.INIT=8'h8E;
  LUT6 un7_0_0_axb_24_cZ(.I0(un7_0_6[23:23]),.I1(un7_0_10[23:23]),.I2(un7_0_6[24:24]),.I3(un7_0_10[24:24]),.I4(un7_0_8[23:23]),.I5(un7_0_8[24:24]),.O(un7_0_0_axb_24));
defparam un7_0_0_axb_24_cZ.INIT=64'h1EE17887E11E8778;
  LUT5 ZFF_X2_15_rep1_RNIMQ9A1(.I0(ZFF_X2_15_rep1),.I1(ZFF_X2_10_rep1),.I2(ZFF_X2_14_rep1),.I3(ZFF_X2[9:9]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_8_axb_20));
defparam ZFF_X2_15_rep1_RNIMQ9A1.INIT=32'h99699699;
  LUT6 un9_axb_9_cZ(.I0(ZFF_Y1[5:5]),.I1(ZFF_Y1[6:6]),.I2(un9_8[11:11]),.I3(un9_8[10:10]),.I4(un9_6[11:11]),.I5(un9_6[10:10]),.O(un9_axb_9));
defparam un9_axb_9_cZ.INIT=64'h3C69C39669C3963C;
  LUT5 desc446(.I0(ZFF_X2_fast[3:3]),.I1(ZFF_X2_2_rep1),.I2(ZFF_X2_fast[8:8]),.I3(ZFF_X2_fast[7:7]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_8_axb_13));
defparam desc446.INIT=32'h96A5695A;
  LUT3 un10_8_o5_15_cZ(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[5:5]),.I2(ZFF_Y2[10:10]),.O(un10_8_o5_15));
defparam un10_8_o5_15_cZ.INIT=8'h8E;
  LUT5 un7_0_6_axb_16_cZ(.I0(ZFF_X1_fast[9:9]),.I1(ZFF_X1_2_rep1),.I2(ZFF_X1_1_rep1),.I3(ZFF_X1_8_rep1),.I4(ZFF_X1_fast[16:16]),.O(un7_0_6_axb_16));
defparam un7_0_6_axb_16_cZ.INIT=32'h69669969;
  LUT6 ZFF_X0_4_rep1_RNI7KFF1(.I0(ZFF_X0_2_rep1),.I1(ZFF_X0_4_rep1),.I2(ZFF_X0_3_rep1),.I3(ZFF_X0_14_rep1),.I4(ZFF_X0_1_rep1),.I5(ZFF_X0[13:13]),.O(un6_0_6_axb_9));
defparam ZFF_X0_4_rep1_RNI7KFF1.INIT=64'h9669669999669669;
  LUT6 ZFF_X2_14_rep1_RNII91F1(.I0(ZFF_X2_14_rep1),.I1(ZFF_X2[10:10]),.I2(ZFF_X2[9:9]),.I3(ZFF_X2[15:15]),.I4(ZFF_X2[12:12]),.I5(ZFF_X2[11:11]),.O(un8_0_6_axb_17));
defparam ZFF_X2_14_rep1_RNII91F1.INIT=64'h36C9C9366C93936C;
  LUT3 un10_8_o5_19_cZ(.I0(ZFF_Y2[14:14]),.I1(ZFF_Y2[11:11]),.I2(ZFF_Y2[9:9]),.O(un10_8_o5_19));
defparam un10_8_o5_19_cZ.INIT=8'hD4;
  LUT5 ZFF_X0_16_rep1_RNISNQV(.I0(ZFF_X0_16_rep1),.I1(ZFF_X0[6:6]),.I2(ZFF_X0[7:7]),.I3(ZFF_X0[9:9]),.I4(ZFF_X0[8:8]),.O(un6_0_6_axb_14));
defparam ZFF_X0_16_rep1_RNISNQV.INIT=32'h87781EE1;
  LUT5 desc447(.I0(ZFF_X2[10:10]),.I1(ZFF_X2[15:15]),.I2(ZFF_X2[12:12]),.I3(ZFF_X2[13:13]),.I4(ZFF_X2[11:11]),.O(un8_0_6_axb_18));
defparam desc447.INIT=32'h24DBDB24;
  LUT5 ZFF_X0_15_rep1_RNI781E2(.I0(ZFF_X0_15_rep1),.I1(ZFF_X0[10:10]),.I2(ZFF_X0[12:12]),.I3(ZFF_X0[11:11]),.I4(ZFF_X0[13:13]),.O(un6_0_6_axb_18));
defparam ZFF_X0_15_rep1_RNI781E2.INIT=32'h42BDBD42;
  LUT6 un6_0_0_axb_21_cZ(.I0(un6_0_8[20:20]),.I1(un6_0_8[21:21]),.I2(un6_0_9[20:20]),.I3(un6_0_9[21:21]),.I4(un6_0_6[20:20]),.I5(un6_0_6[21:21]),.O(un6_0_0_axb_21));
defparam un6_0_0_axb_21_cZ.INIT=64'h36C96C93C936936C;
  LUT2 un7_0_10_o5_21_cZ(.I0(ZFF_X1[14:14]),.I1(ZFF_X1[11:11]),.O(un7_0_10_o5_21));
defparam un7_0_10_o5_21_cZ.INIT=4'hD;
  LUT2 un7_0_10_o5_19_cZ(.I0(ZFF_X1[12:12]),.I1(ZFF_X1[9:9]),.O(un7_0_10_o5_19));
defparam un7_0_10_o5_19_cZ.INIT=4'hD;
  LUT6 ZFF_X2_15_rep1_RNITMOI1(.I0(ZFF_X2_15_rep1),.I1(ZFF_X2_2_rep1),.I2(ZFF_X2[3:3]),.I3(ZFF_X2_14_rep1),.I4(ZFF_X2[4:4]),.I5(ZFF_X2[5:5]),.O(un8_0_6_axb_10));
defparam ZFF_X2_15_rep1_RNITMOI1.INIT=64'h96A55A96695AA569;
  LUT5 ZFF_X0_16_rep1_RNIOJQV(.I0(ZFF_X0_16_rep1),.I1(ZFF_X0[6:6]),.I2(ZFF_X0[7:7]),.I3(ZFF_X0[5:5]),.I4(ZFF_X0[8:8]),.O(un6_0_6_axb_13));
defparam ZFF_X0_16_rep1_RNIOJQV.INIT=32'h93366CC9;
  LUT5 ZFF_X0_6_rep1_RNIGNIT(.I0(ZFF_X0_6_rep1),.I1(ZFF_X0_4_rep1),.I2(ZFF_X0_16_rep1),.I3(ZFF_X0[7:7]),.I4(ZFF_X0[5:5]),.O(un6_0_6_axb_12));
defparam ZFF_X0_6_rep1_RNIGNIT.INIT=32'h817E7E81;
  LUT6 ZFF_Y1_1_rep1_RNILNPM1(.I0(un9_8_6_rep1),.I1(ZFF_Y1_6_rep1),.I2(ZFF_Y1_3_rep1),.I3(ZFF_Y1[4:4]),.I4(ZFF_Y1_7_rep1),.I5(un9_10_8_rep1),.O(un9_10_axb_14));
defparam ZFF_Y1_1_rep1_RNILNPM1.INIT=64'h56A9A9566A95956A;
  LUT3 un10_8_o5_12_cZ(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[2:2]),.O(un10_8_o5_12));
defparam un10_8_o5_12_cZ.INIT=8'hD4;
  LUT5 un10_8_ac0_5_cZ(.I0(ZFF_Y2_fast[14:14]),.I1(ZFF_Y2_fast[8:8]),.I2(ZFF_Y2_fast[7:7]),.I3(ZFF_Y2_fast[6:6]),.I4(ZFF_Y2_fast[17:17]),.O(un10_8_ac0_5));
defparam un10_8_ac0_5_cZ.INIT=32'h00020000;
  LUT5 desc448(.I0(ZFF_X0_fast[4:4]),.I1(ZFF_X0_fast[7:7]),.I2(ZFF_X0_fast[6:6]),.I3(ZFF_X0_fast[8:8]),.I4(ZFF_X0_fast[5:5]),.O(un6_0_8_axb_3));
defparam desc448.INIT=32'h1EE18778;
  LUT5 desc449(.I0(ZFF_X1_fast[10:10]),.I1(ZFF_X1_fast[6:6]),.I2(ZFF_X1_0_rep1),.I3(ZFF_X1_7_rep1),.I4(ZFF_X1_fast[16:16]),.O(un7_0_6_axb_14));
defparam desc449.INIT=32'h7887E11E;
  LUT6 un8_0_0_axb_15_cZ(.I0(ZFF_X2[7:7]),.I1(ZFF_X2[8:8]),.I2(un8_0_8[14:14]),.I3(un8_0_8[15:15]),.I4(un8_0_6[14:14]),.I5(un8_0_6[15:15]),.O(un8_0_0_axb_15));
defparam un8_0_0_axb_15_cZ.INIT=64'h9669669969969966;
  LUT3 un10_8_o5_23_cZ(.I0(ZFF_Y2[13:13]),.I1(ZFF_Y2[15:15]),.I2(ZFF_Y2[17:17]),.O(un10_8_o5_23));
defparam un10_8_o5_23_cZ.INIT=8'h8E;
  LUT6 un8_0_0_axb_17_cZ(.I0(un8_0_8[16:16]),.I1(un8_0_8[17:17]),.I2(un8_0_9[16:16]),.I3(un8_0_9[17:17]),.I4(un8_0_6[16:16]),.I5(un8_0_6[17:17]),.O(un8_0_0_axb_17));
defparam un8_0_0_axb_17_cZ.INIT=64'h36C96C93C936936C;
  LUT6 ZFF_Y1_14_rep1_RNI5G341(.I0(un9_11_26_rep1),.I1(ZFF_Y1_6_rep1),.I2(ZFF_Y1_3_rep1),.I3(ZFF_Y1_5_rep1),.I4(un9_10_8_rep1),.I5(un9_8[7:7]),.O(un9_10_axb_13));
defparam ZFF_Y1_14_rep1_RNI5G341.INIT=64'h3C69C39669C3963C;
  LUT6 desc450(.I0(ZFF_X1_fast[5:5]),.I1(ZFF_X1_3_rep1),.I2(ZFF_X1_fast[2:2]),.I3(ZFF_X1_fast[6:6]),.I4(ZFF_X1_1_rep1),.I5(ZFF_X1_0_rep1),.O(un7_0_8_axb_6));
defparam desc450.INIT=64'h36C9C9366C93936C;
  LUT5 un10_10_cZ(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[5:5]),.I3(ZFF_Y2[3:3]),.I4(ZFF_Y2[1:1]),.O(un10_10));
defparam un10_10_cZ.INIT=32'h00000002;
  LUT6 un8_0_0_axb_23_cZ(.I0(un8_0_8[22:22]),.I1(un8_0_8[23:23]),.I2(un8_0_9[22:22]),.I3(un8_0_9[23:23]),.I4(un8_0_6[22:22]),.I5(un8_0_6[23:23]),.O(un8_0_0_axb_23));
defparam un8_0_0_axb_23_cZ.INIT=64'h36C96C93C936936C;
  LUT5 desc451(.I0(ZFF_X1_fast[12:12]),.I1(ZFF_X1_fast[11:11]),.I2(ZFF_X1_fast[3:3]),.I3(ZFF_X1_fast[2:2]),.I4(ZFF_X1_1_rep1),.O(un7_0_6_axb_9));
defparam desc451.INIT=32'h69965AA5;
  LUT6 ZFF_X1_2_rep1_RNI7F391(.I0(ZFF_X1_2_rep1),.I1(ZFF_X1_12_rep1),.I2(ZFF_X1_3_rep1),.I3(ZFF_X1_11_rep1),.I4(ZFF_X1_10_rep1),.I5(ZFF_X1_13_rep1),.O(un7_0_8_axb_16));
defparam ZFF_X1_2_rep1_RNI7F391.INIT=64'h1EE17887E11E8778;
  LUT6 desc452(.I0(ZFF_X0_fast[13:13]),.I1(ZFF_X0_2_rep1),.I2(ZFF_X0_12_rep1),.I3(ZFF_X0_3_rep1),.I4(ZFF_X0_fast[0:0]),.I5(ZFF_X0_1_rep1),.O(un6_0_6_axb_8));
defparam desc452.INIT=64'h9A6559A6659AA659;
  LUT3 un10_8_o5_21_cZ(.I0(ZFF_Y2[11:11]),.I1(ZFF_Y2[13:13]),.I2(ZFF_Y2[16:16]),.O(un10_8_o5_21));
defparam un10_8_o5_21_cZ.INIT=8'h8E;
  LUT6 desc453(.I0(ZFF_X2_fast[13:13]),.I1(ZFF_X2_2_rep1),.I2(ZFF_X2_3_rep1),.I3(ZFF_X2_fast[1:1]),.I4(ZFF_X2_fast[0:0]),.I5(ZFF_X2_fast[12:12]),.O(un8_0_6_axb_8));
defparam desc453.INIT=64'h96695AA5A55A9669;
  LUT6 ZFF_X0_11_rep1_RNIV6V71(.I0(ZFF_X0_11_rep1),.I1(ZFF_X0_6_rep1),.I2(ZFF_X0_10_rep1),.I3(ZFF_X0_fast[0:0]),.I4(ZFF_X0_1_rep1),.I5(ZFF_X0_fast[5:5]),.O(un6_0_6_axb_6));
defparam ZFF_X0_11_rep1_RNIV6V71.INIT=64'h9969669669669699;
  LUT3 Y_out_double_2_6_0_o5_14_cZ(.I0(pgZFF_X1[14:14]),.I1(pgZFF_Y1[14:14]),.I2(pgZFF_Y2[14:14]),.O(Y_out_double_2_6_0_o5_14));
defparam Y_out_double_2_6_0_o5_14_cZ.INIT=8'h2B;
  LUT4 un6_0_0_o5_15_cZ(.I0(ZFF_X0[7:7]),.I1(ZFF_X0[8:8]),.I2(un6_0_8[15:15]),.I3(un6_0_6[15:15]),.O(un6_0_0_o5_15));
defparam un6_0_0_o5_15_cZ.INIT=16'hF660;
  LUT6 un7_0_0_axb_14_cZ(.I0(ZFF_X1[7:7]),.I1(ZFF_X1[11:11]),.I2(un7_0_6[13:13]),.I3(un7_0_6[14:14]),.I4(un7_0_8[13:13]),.I5(un7_0_8[14:14]),.O(un7_0_0_axb_14));
defparam un7_0_0_axb_14_cZ.INIT=64'h36C96C93C936936C;
  LUT6 desc454(.I0(ZFF_X1_fast[12:12]),.I1(ZFF_X1_4_rep1),.I2(ZFF_X1_fast[5:5]),.I3(ZFF_X1_3_rep1),.I4(ZFF_X1_6_rep1),.I5(ZFF_X1_fast[14:14]),.O(un7_0_8_axb_9));
defparam desc454.INIT=64'h6669999669999666;
  LUT6 ZFF_X2_2_rep1_RNIPS3B1(.I0(ZFF_X2_2_rep1),.I1(ZFF_X2[3:3]),.I2(ZFF_X2_14_rep1),.I3(ZFF_X2[4:4]),.I4(ZFF_X2[1:1]),.I5(ZFF_X2[13:13]),.O(un8_0_6_axb_9));
defparam ZFF_X2_2_rep1_RNIPS3B1.INIT=64'h96695AA5A55A9669;
  LUT2 un7_0_6_o5_20_cZ(.I0(ZFF_X1_13_rep1),.I1(ZFF_X1[6:6]),.O(un7_0_6_o5_20));
defparam un7_0_6_o5_20_cZ.INIT=4'hB;
  LUT6 un7_0_0_axb_21_cZ(.I0(un7_0_6[20:20]),.I1(un7_0_10[20:20]),.I2(un7_0_6[21:21]),.I3(un7_0_10[21:21]),.I4(un7_0_8[20:20]),.I5(un7_0_8[21:21]),.O(un7_0_0_axb_21));
defparam un7_0_0_axb_21_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 desc455(.I0(ZFF_X1_fast[7:7]),.I1(ZFF_X1_4_rep1),.I2(ZFF_X1_3_rep1),.I3(ZFF_X1_fast[2:2]),.I4(ZFF_X1_fast[6:6]),.I5(ZFF_X1_1_rep1),.O(un7_0_8_axb_7));
defparam desc455.INIT=64'h6699699669969966;
  LUT5 ZFF_X2_6_rep1_RNIRAU31(.I0(ZFF_X2_6_rep1),.I1(ZFF_X2_fast[11:11]),.I2(ZFF_X2_10_rep1),.I3(ZFF_X2_fast[5:5]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_8_axb_16));
defparam ZFF_X2_6_rep1_RNIRAU31.INIT=32'h66969699;
  LUT5 ZFF_X0_11_rep1_RNI2CH31(.I0(ZFF_X0_11_rep1),.I1(ZFF_X0_6_rep1),.I2(ZFF_X0_10_rep1),.I3(ZFF_X0_fast[5:5]),.I4(ZFF_X0_fast[16:16]),.O(un6_0_8_axb_16));
defparam ZFF_X0_11_rep1_RNI2CH31.INIT=32'h66969699;
  LUT6 desc456(.I0(un9_11_fast[25:25]),.I1(un9_8_6_rep1),.I2(un9_8_7_rep1),.I3(un9_11_26_rep1),.I4(ZFF_Y1[4:4]),.I5(ZFF_Y1_5_rep1),.O(un9_10_axb_12));
defparam desc456.INIT=64'h1EE17887E11E8778;
  LUT6 ZFF_X2_6_rep1_RNIS89T1(.I0(ZFF_X2_6_rep1),.I1(ZFF_X2_fast[1:1]),.I2(ZFF_X2_10_rep1),.I3(ZFF_X2_fast[0:0]),.I4(ZFF_X2_fast[5:5]),.I5(ZFF_X2[11:11]),.O(un8_0_6_axb_6));
defparam ZFF_X2_6_rep1_RNIS89T1.INIT=64'h9969696666969699;
  LUT5 un10_8_axbxc3(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[7:7]),.I2(ZFF_Y2[6:6]),.I3(ZFF_Y2[14:14]),.I4(ZFF_Y2[17:17]),.O(un10_8[17:17]));
defparam un10_8_axbxc3.INIT=32'hFEFF0100;
  LUT4 un10_8_axbxc2(.I0(ZFF_Y2_fast[14:14]),.I1(ZFF_Y2_fast[7:7]),.I2(ZFF_Y2_6_rep1),.I3(ZFF_Y2_8_rep1),.O(un10_8[16:16]));
defparam un10_8_axbxc2.INIT=16'h02FD;
  LUT6 un7_0_0_axb_29_cZ(.I0(un7_0_6[28:28]),.I1(un7_0_10[28:28]),.I2(un7_0_6[29:29]),.I3(un7_0_10[29:29]),.I4(un7_0_8[28:28]),.I5(un7_0_8[29:29]),.O(un7_0_0_axb_29));
defparam un7_0_0_axb_29_cZ.INIT=64'h1EE17887E11E8778;
  LUT3 un10_o5_13_cZ(.I0(ZFF_Y2[13:13]),.I1(un10_8[19:19]),.I2(un10_6[19:19]),.O(un10_o5_13));
defparam un10_o5_13_cZ.INIT=8'hD4;
  LUT6 un7_0_0_axb_32_cZ(.I0(un7_0_6[31:31]),.I1(un7_0_10[31:31]),.I2(un7_0_6[32:32]),.I3(un7_0_10[32:32]),.I4(un7_0_8[31:31]),.I5(un7_0_8[32:32]),.O(un7_0_0_axb_32));
defparam un7_0_0_axb_32_cZ.INIT=64'h1EE17887E11E8778;
  LUT3 un10_o5_15_cZ(.I0(ZFF_Y2[15:15]),.I1(un10_8[21:21]),.I2(un10_6[21:21]),.O(un10_o5_15));
defparam un10_o5_15_cZ.INIT=8'hD4;
  LUT3 un10_o5_16_cZ(.I0(ZFF_Y2[16:16]),.I1(un10_8[22:22]),.I2(un10_6[22:22]),.O(un10_o5_16));
defparam un10_o5_16_cZ.INIT=8'hD4;
  LUT6 un8_0_0_axb_19_cZ(.I0(un8_0_8[18:18]),.I1(un8_0_8[19:19]),.I2(un8_0_9[18:18]),.I3(un8_0_9[19:19]),.I4(un8_0_6[18:18]),.I5(un8_0_6[19:19]),.O(un8_0_0_axb_19));
defparam un8_0_0_axb_19_cZ.INIT=64'h36C96C93C936936C;
  LUT3 un10_o5_19_cZ(.I0(ZFF_Y2[17:17]),.I1(un10_8[25:25]),.I2(un10_6[25:25]),.O(un10_o5_19));
defparam un10_o5_19_cZ.INIT=8'hD4;
  LUT3 un10_o5_20_cZ(.I0(ZFF_Y2[17:17]),.I1(un10_8[26:26]),.I2(un10_6[26:26]),.O(un10_o5_20));
defparam un10_o5_20_cZ.INIT=8'hD4;
  LUT3 un10_o5_21_cZ(.I0(ZFF_Y2[17:17]),.I1(un10_8[27:27]),.I2(un10_6[27:27]),.O(un10_o5_21));
defparam un10_o5_21_cZ.INIT=8'hD4;
  LUT3 un10_o5_22_cZ(.I0(ZFF_Y2[17:17]),.I1(un10_8[28:28]),.I2(un10_6[28:28]),.O(un10_o5_22));
defparam un10_o5_22_cZ.INIT=8'hD4;
  LUT6 desc457(.I0(ZFF_Y1[9:9]),.I1(un9_11_25_rep1),.I2(un9_11[24:24]),.I3(ZFF_Y1[15:15]),.I4(ZFF_Y1_16_rep1),.I5(un9_11[22:22]),.O(un9_10_axb_23));
defparam desc457.INIT=64'h366CC993C993366C;
  LUT6 un8_0_0_axb_28_cZ(.I0(un8_0_6[28:28]),.I1(un8_0_8[28:28]),.I2(un8_0_8[27:27]),.I3(un8_0_9[28:28]),.I4(un8_0_9[27:27]),.I5(un8_0_6[27:27]),.O(un8_0_0_axb_28));
defparam un8_0_0_axb_28_cZ.INIT=64'h6699699669969966;
  LUT6 desc458(.I0(ZFF_Y1[9:9]),.I1(un9_11_23_rep1),.I2(ZFF_Y1[8:8]),.I3(un9_11[24:24]),.I4(ZFF_Y1[15:15]),.I5(un9_11[26:26]),.O(un9_10_axb_22));
defparam desc458.INIT=64'h56A9A9566A95956A;
  LUT5 desc459(.I0(ZFF_X2[10:10]),.I1(ZFF_X2[9:9]),.I2(ZFF_X2[7:7]),.I3(ZFF_X2[8:8]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_6_axb_15));
defparam desc459.INIT=32'h956A56A9;
  LUT6 ZFF_Y1_11_rep1_RNI14NT1(.I0(ZFF_Y1[7:7]),.I1(un9_11_23_rep1),.I2(un9_11_25_rep1),.I3(ZFF_Y1[8:8]),.I4(un9_11[22:22]),.I5(un9_11[26:26]),.O(un9_10_axb_21));
defparam ZFF_Y1_11_rep1_RNI14NT1.INIT=64'h36C96C93C936936C;
  LUT3 un10_8_o5_11_cZ(.I0(ZFF_Y2[6:6]),.I1(ZFF_Y2[3:3]),.I2(ZFF_Y2[1:1]),.O(un10_8_o5_11));
defparam un10_8_o5_11_cZ.INIT=8'hD4;
  LUT6 ZFF_X1_6_rep1_RNIGKQQ1(.I0(ZFF_X1_6_rep1),.I1(ZFF_X1_9_rep1),.I2(ZFF_X1_7_rep1),.I3(ZFF_X1_15_rep1),.I4(ZFF_X1_fast[14:14]),.I5(ZFF_X1_8_rep1),.O(un7_0_8_axb_12));
defparam ZFF_X1_6_rep1_RNIGKQQ1.INIT=64'h3CC369966996C33C;
  LUT6 ZFF_Y1_11_rep1_RNITJFK1(.I0(ZFF_Y1_6_rep1),.I1(un9_11_23_rep1),.I2(un9_11_24_rep1),.I3(ZFF_Y1_7_rep1),.I4(ZFF_Y1_15_rep1),.I5(ZFF_Y1_16_rep1),.O(un9_6_0_axb_24));
defparam ZFF_Y1_11_rep1_RNITJFK1.INIT=64'h1EE17887E11E8778;
  LUT6 ZFF_Y1_9_rep1_RNI593K1(.I0(ZFF_Y1_9_rep1),.I1(un9_11_23_rep1),.I2(un9_11_24_rep1),.I3(ZFF_Y1[5:5]),.I4(ZFF_Y1[6:6]),.I5(ZFF_Y1[8:8]),.O(un9_10_axb_19));
defparam ZFF_Y1_9_rep1_RNI593K1.INIT=64'h5A69A59669A5965A;
  LUT6 desc460(.I0(ZFF_X1_fast[7:7]),.I1(ZFF_X1_4_rep1),.I2(ZFF_X1_fast[5:5]),.I3(ZFF_X1_3_rep1),.I4(ZFF_X1_fast[2:2]),.I5(ZFF_X1_fast[14:14]),.O(un7_0_8_axb_8));
defparam desc460.INIT=64'h1EE17887E11E8778;
  LUT3 un9_8_o5_13_cZ(.I0(ZFF_Y1_fast[17:17]),.I1(ZFF_Y1_fast[7:7]),.I2(un9_10_8_rep1),.O(un9_8_o5_13));
defparam un9_8_o5_13_cZ.INIT=8'h71;
  LUT3 un9_8_o5_17_cZ(.I0(ZFF_Y1_17_rep1),.I1(un9_11_fast[23:23]),.I2(ZFF_Y1_4_rep1),.O(un9_8_o5_17));
defparam un9_8_o5_17_cZ.INIT=8'h71;
  LUT5 desc461(.I0(ZFF_X0_fast[1:1]),.I1(ZFF_X0_fast[10:10]),.I2(ZFF_X0_fast[11:11]),.I3(ZFF_X0_fast[0:0]),.I4(ZFF_X0_fast[9:9]),.O(un6_0_8_axb_6));
defparam desc461.INIT=32'h96A5695A;
  LUT6 desc462(.I0(un9_11_fast[25:25]),.I1(un9_8_6_rep1),.I2(un9_11_24_rep1),.I3(ZFF_Y1_3_rep1),.I4(ZFF_Y1[4:4]),.I5(un9_10_8_rep1),.O(un9_10_axb_11));
defparam desc462.INIT=64'h6669999669999666;
  LUT6 desc463(.I0(un9_11_fast[25:25]),.I1(un9_8_7_rep1),.I2(un9_11_fast[23:23]),.I3(un9_11_24_rep1),.I4(ZFF_Y1_3_rep1),.I5(un9_10_8_rep1),.O(un9_10_axb_10));
defparam desc463.INIT=64'h17E8E817E81717E8;
  LUT6 desc464(.I0(un9_11_fast[22:22]),.I1(ZFF_Y1_8_rep1),.I2(un9_11_fast[25:25]),.I3(un9_8_6_rep1),.I4(un9_8_7_rep1),.I5(un9_11_fast[23:23]),.O(un9_10_axb_9));
defparam desc464.INIT=64'h1E78E187E1871E78;
  LUT6 un9_axb_15_cZ(.I0(un9_8[16:16]),.I1(un9_8[17:17]),.I2(un9_10[16:16]),.I3(un9_10[17:17]),.I4(un9_6[16:16]),.I5(un9_6[17:17]),.O(un9_axb_15));
defparam un9_axb_15_cZ.INIT=64'h36C96C93C936936C;
  LUT4 un9_o5_10_cZ(.I0(un9_8[7:7]),.I1(un9_10[8:8]),.I2(un9_8[12:12]),.I3(un9_6[12:12]),.O(un9_o5_10));
defparam un9_o5_10_cZ.INIT=16'hF660;
  LUT6 desc465(.I0(un9_11_fast[24:24]),.I1(un9_11_fast[25:25]),.I2(ZFF_Y1_6_rep1),.I3(ZFF_Y1_fast[8:8]),.I4(ZFF_Y1_5_rep1),.I5(ZFF_Y1_7_rep1),.O(un9_10_axb_6));
defparam desc465.INIT=64'h3CC369966996C33C;
  LUT3 un10_8_o5_20_cZ(.I0(ZFF_Y2[12:12]),.I1(ZFF_Y2[10:10]),.I2(ZFF_Y2[15:15]),.O(un10_8_o5_20));
defparam un10_8_o5_20_cZ.INIT=8'h8E;
  LUT6 un9_axb_29_cZ(.I0(un9_8[30:30]),.I1(un9_8[31:31]),.I2(un9_10[30:30]),.I3(un9_10[31:31]),.I4(un9_6[30:30]),.I5(un9_6[31:31]),.O(un9_axb_29));
defparam un9_axb_29_cZ.INIT=64'h36C96C93C936936C;
  LUT6 ZFF_X1_11_rep1_RNIDE5U1(.I0(ZFF_X1_11_rep1),.I1(ZFF_X1_1_rep1),.I2(ZFF_X1_10_rep1),.I3(ZFF_X1_9_rep1),.I4(ZFF_X1_0_rep1),.I5(ZFF_X1_8_rep1),.O(un7_0_8_axb_14));
defparam ZFF_X1_11_rep1_RNIDE5U1.INIT=64'h6699699669969966;
  LUT3 un9_cry_7_RNO_cZ(.I0(ZFF_Y1[6:6]),.I1(ZFF_Y1[3:3]),.I2(un9_10[8:8]),.O(un9_cry_7_RNO));
defparam un9_cry_7_RNO_cZ.INIT=8'h90;
  LUT5 desc466(.I0(ZFF_X2[6:6]),.I1(ZFF_X2[9:9]),.I2(ZFF_X2[7:7]),.I3(ZFF_X2[8:8]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_6_axb_14));
defparam desc466.INIT=32'h963C3C69;
  LUT5 desc467(.I0(ZFF_X2[6:6]),.I1(ZFF_X2[5:5]),.I2(ZFF_X2[7:7]),.I3(ZFF_X2[8:8]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_6_axb_13));
defparam desc467.INIT=32'h956A56A9;
  LUT5 desc468(.I0(un9_11_fast[22:22]),.I1(ZFF_Y1_17_rep1),.I2(un9_11_fast[23:23]),.I3(ZFF_Y1_3_rep1),.I4(ZFF_Y1_4_rep1),.O(un9_8_axb_17));
defparam desc468.INIT=32'h3C96C369;
  LUT6 un7_0_0_o5_18_cZ(.I0(ZFF_X1[8:8]),.I1(ZFF_X1[15:15]),.I2(ZFF_X1[9:9]),.I3(ZFF_X1[11:11]),.I4(un7_0_6[18:18]),.I5(un7_0_8[18:18]),.O(un7_0_0_o5_18));
defparam un7_0_0_o5_18_cZ.INIT=64'hFFFFC396C3960000;
  LUT5 desc469(.I0(ZFF_Y1_fast[17:17]),.I1(un9_11_fast[24:24]),.I2(ZFF_Y1_fast[7:7]),.I3(ZFF_Y1_fast[6:6]),.I4(un9_10_8_rep1),.O(un9_8_axb_13));
defparam desc469.INIT=32'hE1781E87;
  LUT2 un7_0_10_o5_20_cZ(.I0(ZFF_X1[10:10]),.I1(ZFF_X1[13:13]),.O(un7_0_10_o5_20));
defparam un7_0_10_o5_20_cZ.INIT=4'hB;
  LUT6 desc470(.I0(ZFF_Y1_fast[17:17]),.I1(un9_11_fast[26:26]),.I2(ZFF_Y1_fast[5:5]),.I3(un9_11_fast[24:24]),.I4(ZFF_Y1_fast[9:9]),.I5(ZFF_Y1_fast[6:6]),.O(un9_8_axb_12));
defparam desc470.INIT=64'h659AA6599A6559A6;
  LUT6 un9_axb_40_cZ(.I0(un9_10[42:42]),.I1(un9_8[42:42]),.I2(un9_8[41:41]),.I3(un9_10[41:41]),.I4(un9_6[42:42]),.I5(un9_6[41:41]),.O(un9_axb_40));
defparam un9_axb_40_cZ.INIT=64'h6669999669999666;
  LUT6 ZFF_Y1_8_rep1_RNITLG52(.I0(ZFF_Y1_8_rep1),.I1(un9_8_6_rep1),.I2(ZFF_Y1[4:4]),.I3(ZFF_Y1_5_rep1),.I4(ZFF_Y1_7_rep1),.I5(un9_8[7:7]),.O(un9_10_axb_15));
defparam ZFF_Y1_8_rep1_RNITLG52.INIT=64'h56A96A95A956956A;
  LUT5 ZFF_Y2_14_rep1_RNIRMDL(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2[10:10]),.I2(ZFF_Y2[11:11]),.I3(ZFF_Y2[16:16]),.I4(ZFF_Y2[15:15]),.O(un10_6_axb_20));
defparam ZFF_Y2_14_rep1_RNIRMDL.INIT=32'h2DB4D24B;
  LUT2 un9_8_o5_18_cZ(.I0(un9_11_fast[24:24]),.I1(ZFF_Y1_5_rep1),.O(un9_8_o5_18));
defparam un9_8_o5_18_cZ.INIT=4'hD;
  LUT3 un6_0_8_o5_10_cZ(.I0(ZFF_X0_fast[15:15]),.I1(ZFF_X0_fast[0:0]),.I2(ZFF_X0_fast[5:5]),.O(un6_0_8_o5_10));
defparam un6_0_8_o5_10_cZ.INIT=8'h8E;
  LUT3 Y_out_double_2_6_0_o5_1_cZ(.I0(pgZFF_X1[1:1]),.I1(pgZFF_Y1[1:1]),.I2(pgZFF_Y2[1:1]),.O(Y_out_double_2_6_0_o5_1));
defparam Y_out_double_2_6_0_o5_1_cZ.INIT=8'h2B;
  LUT3 Y_out_double_2_6_0_o5_3_cZ(.I0(pgZFF_X1[3:3]),.I1(pgZFF_Y1[3:3]),.I2(pgZFF_Y2[3:3]),.O(Y_out_double_2_6_0_o5_3));
defparam Y_out_double_2_6_0_o5_3_cZ.INIT=8'h2B;
  LUT3 Y_out_double_2_6_0_o5_5_cZ(.I0(pgZFF_X1[5:5]),.I1(pgZFF_Y1[5:5]),.I2(pgZFF_Y2[5:5]),.O(Y_out_double_2_6_0_o5_5));
defparam Y_out_double_2_6_0_o5_5_cZ.INIT=8'h2B;
  LUT3 Y_out_double_2_6_0_o5_7_cZ(.I0(pgZFF_X1[7:7]),.I1(pgZFF_Y1[7:7]),.I2(pgZFF_Y2[7:7]),.O(Y_out_double_2_6_0_o5_7));
defparam Y_out_double_2_6_0_o5_7_cZ.INIT=8'h2B;
  LUT2 un9_8_s_30(.I0(ZFF_Y1[16:16]),.I1(un9_8_cry_29),.O(un9_8[38:38]));
defparam un9_8_s_30.INIT=4'h9;
  LUT3 Y_out_double_2_6_0_o5_9_cZ(.I0(pgZFF_X1[9:9]),.I1(pgZFF_Y1[9:9]),.I2(pgZFF_Y2[9:9]),.O(Y_out_double_2_6_0_o5_9));
defparam Y_out_double_2_6_0_o5_9_cZ.INIT=8'h2B;
  LUT3 Y_out_double_2_6_0_o5_10_cZ(.I0(pgZFF_X1[10:10]),.I1(pgZFF_Y1[10:10]),.I2(pgZFF_Y2[10:10]),.O(Y_out_double_2_6_0_o5_10));
defparam Y_out_double_2_6_0_o5_10_cZ.INIT=8'h2B;
  LUT3 Y_out_double_2_6_0_o5_11_cZ(.I0(pgZFF_X1[11:11]),.I1(pgZFF_Y1[11:11]),.I2(pgZFF_Y2[11:11]),.O(Y_out_double_2_6_0_o5_11));
defparam Y_out_double_2_6_0_o5_11_cZ.INIT=8'h2B;
  LUT3 Y_out_double_2_6_0_o5_13_cZ(.I0(pgZFF_X1[13:13]),.I1(pgZFF_Y1[13:13]),.I2(pgZFF_Y2[13:13]),.O(Y_out_double_2_6_0_o5_13));
defparam Y_out_double_2_6_0_o5_13_cZ.INIT=8'h2B;
  LUT6 un8_0_0_axb_21_cZ(.I0(un8_0_8[20:20]),.I1(un8_0_8[21:21]),.I2(un8_0_9[20:20]),.I3(un8_0_9[21:21]),.I4(un8_0_6[20:20]),.I5(un8_0_6[21:21]),.O(un8_0_0_axb_21));
defparam un8_0_0_axb_21_cZ.INIT=64'h36C96C93C936936C;
  LUT3 Y_out_double_2_6_0_o5_15_cZ(.I0(pgZFF_X1[15:15]),.I1(pgZFF_Y1[15:15]),.I2(pgZFF_Y2[15:15]),.O(Y_out_double_2_6_0_o5_15));
defparam Y_out_double_2_6_0_o5_15_cZ.INIT=8'h2B;
  LUT6 un8_0_0_axb_24_cZ(.I0(un8_0_8[23:23]),.I1(un8_0_8[24:24]),.I2(un8_0_9[23:23]),.I3(un8_0_9[24:24]),.I4(un8_0_6[23:23]),.I5(un8_0_6[24:24]),.O(un8_0_0_axb_24));
defparam un8_0_0_axb_24_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un8_0_0_axb_25_cZ(.I0(un8_0_8[24:24]),.I1(un8_0_8[25:25]),.I2(un8_0_9[24:24]),.I3(un8_0_9[25:25]),.I4(un8_0_6[24:24]),.I5(un8_0_6[25:25]),.O(un8_0_0_axb_25));
defparam un8_0_0_axb_25_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un8_0_0_axb_26_cZ(.I0(un8_0_8[25:25]),.I1(un8_0_8[26:26]),.I2(un8_0_9[25:25]),.I3(un8_0_9[26:26]),.I4(un8_0_6[25:25]),.I5(un8_0_6[26:26]),.O(un8_0_0_axb_26));
defparam un8_0_0_axb_26_cZ.INIT=64'h36C96C93C936936C;
  LUT6 ZFF_X1_2_rep1_RNIQEKB1(.I0(ZFF_X1_2_rep1),.I1(ZFF_X1_12_rep1),.I2(ZFF_X1_11_rep1),.I3(ZFF_X1_1_rep1),.I4(ZFF_X1_10_rep1),.I5(ZFF_X1_9_rep1),.O(un7_0_8_axb_15));
defparam ZFF_X1_2_rep1_RNIQEKB1.INIT=64'h6669999669999666;
  LUT5 un6_0_0_axb_37_cZ(.I0(ZFF_X0[16:16]),.I1(un6_0_8[36:36]),.I2(un6_0_8[37:37]),.I3(un6_0_9[36:36]),.I4(un6_0_9[37:37]),.O(un6_0_0_axb_37));
defparam un6_0_0_axb_37_cZ.INIT=32'h5A69A596;
  LUT6 ZFF_X1_10_rep1_RNIN0BL1(.I0(ZFF_X1_10_rep1),.I1(ZFF_X1_9_rep1),.I2(ZFF_X1_0_rep1),.I3(ZFF_X1_7_rep1),.I4(ZFF_X1_15_rep1),.I5(ZFF_X1_8_rep1),.O(un7_0_8_axb_13));
defparam ZFF_X1_10_rep1_RNIN0BL1.INIT=64'h5A6969A5A596965A;
  LUT6 ZFF_X0_4_rep1_RNIN2HE1(.I0(ZFF_X0_2_rep1),.I1(ZFF_X0_4_rep1),.I2(ZFF_X0_10_rep1),.I3(ZFF_X0_fast[0:0]),.I4(ZFF_X0_fast[5:5]),.I5(ZFF_X0[9:9]),.O(un6_0_6_axb_5));
defparam ZFF_X0_4_rep1_RNIN2HE1.INIT=64'h87787887E11E1EE1;
  LUT4 un7_0_0_o5_17_cZ(.I0(ZFF_X1[8:8]),.I1(ZFF_X1[11:11]),.I2(un7_0_6[17:17]),.I3(un7_0_8[17:17]),.O(un7_0_0_o5_17));
defparam un7_0_0_o5_17_cZ.INIT=16'hF990;
  LUT6 ZFF_Y1_8_rep1_RNI18OT1(.I0(ZFF_Y1_8_rep1),.I1(un9_11_24_rep1),.I2(un9_11_25_rep1),.I3(ZFF_Y1_7_rep1),.I4(ZFF_Y1_15_rep1),.I5(ZFF_Y1_16_rep1),.O(un9_6_0_axb_25));
defparam ZFF_Y1_8_rep1_RNI18OT1.INIT=64'h5A69A59669A5965A;
  LUT6 un7_0_0_axb_12_cZ(.I0(ZFF_X1[2:2]),.I1(ZFF_X1[6:6]),.I2(un7_0_6[11:11]),.I3(un7_0_6[12:12]),.I4(un7_0_8[11:11]),.I5(un7_0_8[12:12]),.O(un7_0_0_axb_12));
defparam un7_0_0_axb_12_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un7_0_0_axb_25_cZ(.I0(un7_0_6[24:24]),.I1(un7_0_10[24:24]),.I2(un7_0_6[25:25]),.I3(un7_0_10[25:25]),.I4(un7_0_8[24:24]),.I5(un7_0_8[25:25]),.O(un7_0_0_axb_25));
defparam un7_0_0_axb_25_cZ.INIT=64'h1EE17887E11E8778;
  LUT3 Y_out_double_2_6_0_o5_4_cZ(.I0(pgZFF_X1[4:4]),.I1(pgZFF_Y1[4:4]),.I2(pgZFF_Y2[4:4]),.O(Y_out_double_2_6_0_o5_4));
defparam Y_out_double_2_6_0_o5_4_cZ.INIT=8'h2B;
  LUT6 un7_0_0_axb_30_cZ(.I0(un7_0_6[29:29]),.I1(un7_0_10[29:29]),.I2(un7_0_6[30:30]),.I3(un7_0_10[30:30]),.I4(un7_0_8[29:29]),.I5(un7_0_8[30:30]),.O(un7_0_0_axb_30));
defparam un7_0_0_axb_30_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 un7_0_0_axb_31_cZ(.I0(un7_0_6[30:30]),.I1(un7_0_10[30:30]),.I2(un7_0_6[31:31]),.I3(un7_0_10[31:31]),.I4(un7_0_8[30:30]),.I5(un7_0_8[31:31]),.O(un7_0_0_axb_31));
defparam un7_0_0_axb_31_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 un9_axb_14_cZ(.I0(un9_8[15:15]),.I1(un9_8[16:16]),.I2(un9_10[15:15]),.I3(un9_10[16:16]),.I4(un9_6[15:15]),.I5(un9_6[16:16]),.O(un9_axb_14));
defparam un9_axb_14_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un7_0_0_axb_33_cZ(.I0(un7_0_6[33:33]),.I1(un7_0_10[33:33]),.I2(un7_0_6[32:32]),.I3(un7_0_10[32:32]),.I4(un7_0_8[33:33]),.I5(un7_0_8[32:32]),.O(un7_0_0_axb_33));
defparam un7_0_0_axb_33_cZ.INIT=64'h6669999669999666;
  LUT6 un6_0_0_axb_18_cZ(.I0(un6_0_8[17:17]),.I1(un6_0_8[18:18]),.I2(un6_0_9[17:17]),.I3(un6_0_9[18:18]),.I4(un6_0_6[17:17]),.I5(un6_0_6[18:18]),.O(un6_0_0_axb_18));
defparam un6_0_0_axb_18_cZ.INIT=64'h36C96C93C936936C;
  LUT3 un10_o5_17_cZ(.I0(ZFF_Y2[15:15]),.I1(un10_8[23:23]),.I2(un10_6[23:23]),.O(un10_o5_17));
defparam un10_o5_17_cZ.INIT=8'hD4;
  LUT3 un10_o5_18_cZ(.I0(ZFF_Y2[16:16]),.I1(un10_8[24:24]),.I2(un10_6[24:24]),.O(un10_o5_18));
defparam un10_o5_18_cZ.INIT=8'hD4;
  LUT6 un9_axb_19_cZ(.I0(un9_8[20:20]),.I1(un9_8[21:21]),.I2(un9_10[20:20]),.I3(un9_10[21:21]),.I4(un9_6[20:20]),.I5(un9_6[21:21]),.O(un9_axb_19));
defparam un9_axb_19_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_22_cZ(.I0(un6_0_8[21:21]),.I1(un6_0_8[22:22]),.I2(un6_0_9[21:21]),.I3(un6_0_9[22:22]),.I4(un6_0_6[21:21]),.I5(un6_0_6[22:22]),.O(un6_0_0_axb_22));
defparam un6_0_0_axb_22_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_23_cZ(.I0(un6_0_8[22:22]),.I1(un6_0_8[23:23]),.I2(un6_0_9[22:22]),.I3(un6_0_9[23:23]),.I4(un6_0_6[22:22]),.I5(un6_0_6[23:23]),.O(un6_0_0_axb_23));
defparam un6_0_0_axb_23_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_24_cZ(.I0(un6_0_8[23:23]),.I1(un6_0_8[24:24]),.I2(un6_0_9[23:23]),.I3(un6_0_9[24:24]),.I4(un6_0_6[23:23]),.I5(un6_0_6[24:24]),.O(un6_0_0_axb_24));
defparam un6_0_0_axb_24_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_25_cZ(.I0(un6_0_8[24:24]),.I1(un6_0_8[25:25]),.I2(un6_0_9[24:24]),.I3(un6_0_9[25:25]),.I4(un6_0_6[24:24]),.I5(un6_0_6[25:25]),.O(un6_0_0_axb_25));
defparam un6_0_0_axb_25_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_26_cZ(.I0(un6_0_8[25:25]),.I1(un6_0_8[26:26]),.I2(un6_0_9[25:25]),.I3(un6_0_9[26:26]),.I4(un6_0_6[25:25]),.I5(un6_0_6[26:26]),.O(un6_0_0_axb_26));
defparam un6_0_0_axb_26_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_27_cZ(.I0(un6_0_8[26:26]),.I1(un6_0_8[27:27]),.I2(un6_0_9[26:26]),.I3(un6_0_9[27:27]),.I4(un6_0_6[26:26]),.I5(un6_0_6[27:27]),.O(un6_0_0_axb_27));
defparam un6_0_0_axb_27_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_28_cZ(.I0(un6_0_6[28:28]),.I1(un6_0_8[28:28]),.I2(un6_0_8[27:27]),.I3(un6_0_9[28:28]),.I4(un6_0_9[27:27]),.I5(un6_0_6[27:27]),.O(un6_0_0_axb_28));
defparam un6_0_0_axb_28_cZ.INIT=64'h6699699669969966;
  LUT6 un9_axb_27_cZ(.I0(un9_8[28:28]),.I1(un9_8[29:29]),.I2(un9_10[28:28]),.I3(un9_10[29:29]),.I4(un9_6[28:28]),.I5(un9_6[29:29]),.O(un9_axb_27));
defparam un9_axb_27_cZ.INIT=64'h36C96C93C936936C;
  LUT5 un6_0_0_axb_38_cZ(.I0(ZFF_X0[16:16]),.I1(un6_0_8[37:37]),.I2(un6_0_9[37:37]),.I3(un6_0_9[38:38]),.I4(un6_0_8[38:38]),.O(un6_0_0_axb_38));
defparam un6_0_0_axb_38_cZ.INIT=32'hBD4242BD;
  LUT3 un10_8_o5_22_cZ(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2[12:12]),.I2(ZFF_Y2[17:17]),.O(un10_8_o5_22));
defparam un10_8_o5_22_cZ.INIT=8'h8E;
  LUT6 ZFF_Y1_8_rep1_RNI5S071(.I0(ZFF_Y1_8_rep1),.I1(ZFF_Y1_9_rep1),.I2(un9_11_26_rep1),.I3(un9_11_25_rep1),.I4(ZFF_Y1_15_rep1),.I5(ZFF_Y1_16_rep1),.O(un9_6_0_axb_26));
defparam ZFF_Y1_8_rep1_RNI5S071.INIT=64'h3C6969C3C396963C;
  LUT6 ZFF_Y1_9_rep1_RNII2N52(.I0(ZFF_Y1_9_rep1),.I1(un9_11_24_rep1),.I2(ZFF_Y1[6:6]),.I3(ZFF_Y1_7_rep1),.I4(un9_11[25:25]),.I5(un9_11[22:22]),.O(un9_10_axb_20));
defparam ZFF_Y1_9_rep1_RNII2N52.INIT=64'h17E8E817E81717E8;
  LUT3 un10_8_axbxc1(.I0(ZFF_Y2_fast[14:14]),.I1(ZFF_Y2_fast[6:6]),.I2(ZFF_Y2_7_rep1),.O(un10_8[15:15]));
defparam un10_8_axbxc1.INIT=8'h2D;
  LUT5 un7_0_10_axb_15_cZ(.I0(ZFF_X1[5:5]),.I1(ZFF_X1[8:8]),.I2(ZFF_X1_fast[16:16]),.I3(ZFF_X1[4:4]),.I4(ZFF_X1[7:7]),.O(un7_0_10_axb_15));
defparam un7_0_10_axb_15_cZ.INIT=32'h96669996;
  LUT6 un8_0_0_axb_27_cZ(.I0(un8_0_8[26:26]),.I1(un8_0_8[27:27]),.I2(un8_0_9[26:26]),.I3(un8_0_9[27:27]),.I4(un8_0_6[26:26]),.I5(un8_0_6[27:27]),.O(un8_0_0_axb_27));
defparam un8_0_0_axb_27_cZ.INIT=64'h36C96C93C936936C;
  LUT6 desc471(.I0(ZFF_Y1_fast[16:16]),.I1(ZFF_Y1_fast[15:15]),.I2(ZFF_Y1_fast[3:3]),.I3(ZFF_Y1_fast[4:4]),.I4(un9_11_fast[22:22]),.I5(ZFF_Y1_fast[9:9]),.O(un9_8_axb_10));
defparam desc471.INIT=64'h956A6A95A95656A9;
  LUT5 desc472(.I0(un9_8_fast[6:6]),.I1(ZFF_Y1_fast[5:5]),.I2(un9_11_fast[25:25]),.I3(ZFF_Y1_fast[6:6]),.I4(un9_10_8_rep1),.O(un9_8_axb_7));
defparam desc472.INIT=32'h69966969;
  LUT6 un9_axb_21_cZ(.I0(un9_8[22:22]),.I1(un9_8[23:23]),.I2(un9_10[22:22]),.I3(un9_10[23:23]),.I4(un9_6[22:22]),.I5(un9_6[23:23]),.O(un9_axb_21));
defparam un9_axb_21_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un7_0_0_axb_28_cZ(.I0(un7_0_6[27:27]),.I1(un7_0_10[27:27]),.I2(un7_0_6[28:28]),.I3(un7_0_10[28:28]),.I4(un7_0_8[27:27]),.I5(un7_0_8[28:28]),.O(un7_0_0_axb_28));
defparam un7_0_0_axb_28_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 un9_axb_12_cZ(.I0(un9_8[13:13]),.I1(un9_8[14:14]),.I2(un9_10[13:13]),.I3(un9_10[14:14]),.I4(un9_6[13:13]),.I5(un9_6[14:14]),.O(un9_axb_12));
defparam un9_axb_12_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_13_cZ(.I0(un9_8[14:14]),.I1(un9_8[15:15]),.I2(un9_10[14:14]),.I3(un9_10[15:15]),.I4(un9_6[14:14]),.I5(un9_6[15:15]),.O(un9_axb_13));
defparam un9_axb_13_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_16_cZ(.I0(un9_8[17:17]),.I1(un9_8[18:18]),.I2(un9_10[17:17]),.I3(un9_10[18:18]),.I4(un9_6[17:17]),.I5(un9_6[18:18]),.O(un9_axb_16));
defparam un9_axb_16_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_17_cZ(.I0(un9_8[18:18]),.I1(un9_8[19:19]),.I2(un9_10[18:18]),.I3(un9_10[19:19]),.I4(un9_6[18:18]),.I5(un9_6[19:19]),.O(un9_axb_17));
defparam un9_axb_17_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_18_cZ(.I0(un9_8[19:19]),.I1(un9_8[20:20]),.I2(un9_10[19:19]),.I3(un9_10[20:20]),.I4(un9_6[19:19]),.I5(un9_6[20:20]),.O(un9_axb_18));
defparam un9_axb_18_cZ.INIT=64'h36C96C93C936936C;
  LUT3 Y_out_double_2_6_0_o5_12_cZ(.I0(pgZFF_X1[12:12]),.I1(pgZFF_Y1[12:12]),.I2(pgZFF_Y2[12:12]),.O(Y_out_double_2_6_0_o5_12));
defparam Y_out_double_2_6_0_o5_12_cZ.INIT=8'h2B;
  LUT6 un9_axb_20_cZ(.I0(un9_8[21:21]),.I1(un9_8[22:22]),.I2(un9_10[21:21]),.I3(un9_10[22:22]),.I4(un9_6[21:21]),.I5(un9_6[22:22]),.O(un9_axb_20));
defparam un9_axb_20_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_34_cZ(.I0(un9_8[35:35]),.I1(un9_8[36:36]),.I2(un9_10[35:35]),.I3(un9_10[36:36]),.I4(un9_6[35:35]),.I5(un9_6[36:36]),.O(un9_axb_34));
defparam un9_axb_34_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_22_cZ(.I0(un9_8[23:23]),.I1(un9_8[24:24]),.I2(un9_10[23:23]),.I3(un9_10[24:24]),.I4(un9_6[23:23]),.I5(un9_6[24:24]),.O(un9_axb_22));
defparam un9_axb_22_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_23_cZ(.I0(un9_8[24:24]),.I1(un9_8[25:25]),.I2(un9_10[24:24]),.I3(un9_10[25:25]),.I4(un9_6[24:24]),.I5(un9_6[25:25]),.O(un9_axb_23));
defparam un9_axb_23_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_24_cZ(.I0(un9_8[25:25]),.I1(un9_8[26:26]),.I2(un9_10[25:25]),.I3(un9_10[26:26]),.I4(un9_6[25:25]),.I5(un9_6[26:26]),.O(un9_axb_24));
defparam un9_axb_24_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_25_cZ(.I0(un9_8[26:26]),.I1(un9_8[27:27]),.I2(un9_10[26:26]),.I3(un9_10[27:27]),.I4(un9_6[26:26]),.I5(un9_6[27:27]),.O(un9_axb_25));
defparam un9_axb_25_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_26_cZ(.I0(un9_8[27:27]),.I1(un9_8[28:28]),.I2(un9_10[27:27]),.I3(un9_10[28:28]),.I4(un9_6[27:27]),.I5(un9_6[28:28]),.O(un9_axb_26));
defparam un9_axb_26_cZ.INIT=64'h36C96C93C936936C;
  LUT3 Y_out_double_2_6_0_o5_6_cZ(.I0(pgZFF_X1[6:6]),.I1(pgZFF_Y1[6:6]),.I2(pgZFF_Y2[6:6]),.O(Y_out_double_2_6_0_o5_6));
defparam Y_out_double_2_6_0_o5_6_cZ.INIT=8'h2B;
  LUT6 un9_axb_28_cZ(.I0(un9_8[29:29]),.I1(un9_8[30:30]),.I2(un9_10[29:29]),.I3(un9_10[30:30]),.I4(un9_6[29:29]),.I5(un9_6[30:30]),.O(un9_axb_28));
defparam un9_axb_28_cZ.INIT=64'h36C96C93C936936C;
  LUT4 un9_6_0_cry_27_RNO_cZ(.I0(ZFF_Y1[15:15]),.I1(un9_11[22:22]),.I2(ZFF_Y1[17:17]),.I3(un9_10[8:8]),.O(un9_6_0_cry_27_RNO));
defparam un9_6_0_cry_27_RNO_cZ.INIT=16'h6996;
  LUT6 un9_axb_30_cZ(.I0(un9_8[31:31]),.I1(un9_8[32:32]),.I2(un9_10[31:31]),.I3(un9_10[32:32]),.I4(un9_6[31:31]),.I5(un9_6[32:32]),.O(un9_axb_30));
defparam un9_axb_30_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_31_cZ(.I0(un9_8[32:32]),.I1(un9_8[33:33]),.I2(un9_10[32:32]),.I3(un9_10[33:33]),.I4(un9_6[32:32]),.I5(un9_6[33:33]),.O(un9_axb_31));
defparam un9_axb_31_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_32_cZ(.I0(un9_8[33:33]),.I1(un9_8[34:34]),.I2(un9_10[33:33]),.I3(un9_10[34:34]),.I4(un9_6[33:33]),.I5(un9_6[34:34]),.O(un9_axb_32));
defparam un9_axb_32_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_33_cZ(.I0(un9_8[34:34]),.I1(un9_8[35:35]),.I2(un9_10[34:34]),.I3(un9_10[35:35]),.I4(un9_6[34:34]),.I5(un9_6[35:35]),.O(un9_axb_33));
defparam un9_axb_33_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_35_cZ(.I0(un9_8[36:36]),.I1(un9_8[37:37]),.I2(un9_10[36:36]),.I3(un9_10[37:37]),.I4(un9_6[36:36]),.I5(un9_6[37:37]),.O(un9_axb_35));
defparam un9_axb_35_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un7_0_0_axb_13_cZ(.I0(ZFF_X1[6:6]),.I1(ZFF_X1[7:7]),.I2(un7_0_6[12:12]),.I3(un7_0_6[13:13]),.I4(un7_0_8[12:12]),.I5(un7_0_8[13:13]),.O(un7_0_0_axb_13));
defparam un7_0_0_axb_13_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_38_cZ(.I0(un9_8[39:39]),.I1(un9_8[40:40]),.I2(un9_10[39:39]),.I3(un9_10[40:40]),.I4(un9_6[39:39]),.I5(un9_6[40:40]),.O(un9_axb_38));
defparam un9_axb_38_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un9_axb_39_cZ(.I0(un9_8[40:40]),.I1(un9_8[41:41]),.I2(un9_10[40:40]),.I3(un9_10[41:41]),.I4(un9_6[40:40]),.I5(un9_6[41:41]),.O(un9_axb_39));
defparam un9_axb_39_cZ.INIT=64'h36C96C93C936936C;
  LUT6 desc473(.I0(ZFF_Y2_fast[7:7]),.I1(ZFF_Y2_fast[6:6]),.I2(ZFF_Y2[4:4]),.I3(ZFF_Y2[5:5]),.I4(ZFF_Y2[0:0]),.I5(ZFF_Y2[1:1]),.O(un10_6_axb_10));
defparam desc473.INIT=64'h9A6559A6659AA659;
  LUT5 un9_6_0_axb_21_cZ(.I0(ZFF_Y1_9_rep1),.I1(ZFF_Y1[4:4]),.I2(ZFF_Y1_15_rep1),.I3(ZFF_Y1_16_rep1),.I4(ZFF_Y1[3:3]),.O(un9_6_0_axb_21));
defparam un9_6_0_axb_21_cZ.INIT=32'h69969966;
  LUT6 desc474(.I0(ZFF_Y1_fast[15:15]),.I1(un9_11_fast[26:26]),.I2(ZFF_Y1_fast[3:3]),.I3(un9_8_fast[7:7]),.I4(ZFF_Y1_fast[9:9]),.I5(ZFF_Y1_fast[6:6]),.O(un9_8_axb_9));
defparam desc474.INIT=64'h965A69A5A5965A69;
  LUT2 un9_8_o5_19_cZ(.I0(ZFF_Y1_6_rep1),.I1(un9_11_25_rep1),.O(un9_8_o5_19));
defparam un9_8_o5_19_cZ.INIT=4'hB;
  LUT6 un7_0_0_axb_23_cZ(.I0(un7_0_6[22:22]),.I1(un7_0_10[22:22]),.I2(un7_0_6[23:23]),.I3(un7_0_10[23:23]),.I4(un7_0_8[22:22]),.I5(un7_0_8[23:23]),.O(un7_0_0_axb_23));
defparam un7_0_0_axb_23_cZ.INIT=64'h1EE17887E11E8778;
  LUT3 Y_out_double_2_6_0_o5_2_cZ(.I0(pgZFF_X1[2:2]),.I1(pgZFF_Y1[2:2]),.I2(pgZFF_Y2[2:2]),.O(Y_out_double_2_6_0_o5_2));
defparam Y_out_double_2_6_0_o5_2_cZ.INIT=8'h2B;
  LUT6 un7_0_0_axb_27_cZ(.I0(un7_0_6[26:26]),.I1(un7_0_10[26:26]),.I2(un7_0_6[27:27]),.I3(un7_0_10[27:27]),.I4(un7_0_8[26:26]),.I5(un7_0_8[27:27]),.O(un7_0_0_axb_27));
defparam un7_0_0_axb_27_cZ.INIT=64'h1EE17887E11E8778;
  LUT3 Y_out_double_2_6_0_o5_8_cZ(.I0(pgZFF_X1[8:8]),.I1(pgZFF_Y1[8:8]),.I2(pgZFF_Y2[8:8]),.O(Y_out_double_2_6_0_o5_8));
defparam Y_out_double_2_6_0_o5_8_cZ.INIT=8'h2B;
  LUT2 un9_6_0_s_9(.I0(ZFF_Y1[9:9]),.I1(un9_6_0_cry_8),.O(un9_6[9:9]));
defparam un9_6_0_s_9.INIT=4'h9;
  LUT6 un6_0_0_axb_20_cZ(.I0(un6_0_8[19:19]),.I1(un6_0_8[20:20]),.I2(un6_0_9[19:19]),.I3(un6_0_9[20:20]),.I4(un6_0_6[19:19]),.I5(un6_0_6[20:20]),.O(un6_0_0_axb_20));
defparam un6_0_0_axb_20_cZ.INIT=64'h36C96C93C936936C;
  LUT5 ZFF_Y2_6_rep1_RNI2A1O1(.I0(ZFF_Y2_6_rep1),.I1(ZFF_Y2[0:0]),.I2(ZFF_Y2[3:3]),.I3(ZFF_Y2[2:2]),.I4(ZFF_Y2[1:1]),.O(un10_8_axb_11));
defparam ZFF_Y2_6_rep1_RNI2A1O1.INIT=32'h965A69A5;
  LUT6 un7_0_0_axb_11_cZ(.I0(ZFF_X1[1:1]),.I1(ZFF_X1[2:2]),.I2(un7_0_6[10:10]),.I3(un7_0_6[11:11]),.I4(un7_0_8[10:10]),.I5(un7_0_8[11:11]),.O(un7_0_0_axb_11));
defparam un7_0_0_axb_11_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un8_0_0_axb_22_cZ(.I0(un8_0_8[21:21]),.I1(un8_0_8[22:22]),.I2(un8_0_9[21:21]),.I3(un8_0_9[22:22]),.I4(un8_0_6[21:21]),.I5(un8_0_6[22:22]),.O(un8_0_0_axb_22));
defparam un8_0_0_axb_22_cZ.INIT=64'h36C96C93C936936C;
  LUT4 un8_0_0_o5_15_cZ(.I0(ZFF_X2[7:7]),.I1(ZFF_X2[8:8]),.I2(un8_0_8[15:15]),.I3(un8_0_6[15:15]),.O(un8_0_0_o5_15));
defparam un8_0_0_o5_15_cZ.INIT=16'hF660;
  LUT5 un8_0_0_axb_37_cZ(.I0(ZFF_X2[16:16]),.I1(un8_0_8[36:36]),.I2(un8_0_8[37:37]),.I3(un8_0_9[36:36]),.I4(un8_0_9[37:37]),.O(un8_0_0_axb_37));
defparam un8_0_0_axb_37_cZ.INIT=32'h5A69A596;
  LUT5 un6_0_8_axb_5_cZ(.I0(ZFF_X0_fast[10:10]),.I1(ZFF_X0_7_rep1),.I2(ZFF_X0_fast[6:6]),.I3(ZFF_X0_fast[0:0]),.I4(ZFF_X0_fast[9:9]),.O(un6_0_8_axb_5));
defparam un6_0_8_axb_5_cZ.INIT=32'hA956956A;
  LUT6 desc475(.I0(ZFF_Y2[4:4]),.I1(ZFF_Y2[3:3]),.I2(ZFF_Y2[2:2]),.I3(ZFF_Y2[1:1]),.I4(ZFF_Y2[16:16]),.I5(ZFF_Y2[15:15]),.O(un10_6_axb_7));
defparam desc475.INIT=64'h96A5695A5A96A569;
  LUT6 un8_0_0_axb_18_cZ(.I0(un8_0_8[17:17]),.I1(un8_0_8[18:18]),.I2(un8_0_9[17:17]),.I3(un8_0_9[18:18]),.I4(un8_0_6[17:17]),.I5(un8_0_6[18:18]),.O(un8_0_0_axb_18));
defparam un8_0_0_axb_18_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un7_0_0_axb_22_cZ(.I0(un7_0_6[21:21]),.I1(un7_0_10[21:21]),.I2(un7_0_6[22:22]),.I3(un7_0_10[22:22]),.I4(un7_0_8[21:21]),.I5(un7_0_8[22:22]),.O(un7_0_0_axb_22));
defparam un7_0_0_axb_22_cZ.INIT=64'h1EE17887E11E8778;
  LUT5 un8_0_0_axb_38_cZ(.I0(ZFF_X2[16:16]),.I1(un8_0_8[37:37]),.I2(un8_0_9[37:37]),.I3(un8_0_9[38:38]),.I4(un8_0_8[38:38]),.O(un8_0_0_axb_38));
defparam un8_0_0_axb_38_cZ.INIT=32'hBD4242BD;
  LUT6 un7_0_0_axb_20_cZ(.I0(un7_0_6[19:19]),.I1(un7_0_10[19:19]),.I2(un7_0_6[20:20]),.I3(un7_0_10[20:20]),.I4(un7_0_8[19:19]),.I5(un7_0_8[20:20]),.O(un7_0_0_axb_20));
defparam un7_0_0_axb_20_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 un7_0_0_axb_26_cZ(.I0(un7_0_6[25:25]),.I1(un7_0_10[25:25]),.I2(un7_0_6[26:26]),.I3(un7_0_10[26:26]),.I4(un7_0_8[25:25]),.I5(un7_0_8[26:26]),.O(un7_0_0_axb_26));
defparam un7_0_0_axb_26_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 desc476(.I0(ZFF_Y2[4:4]),.I1(ZFF_Y2[5:5]),.I2(ZFF_Y2[3:3]),.I3(ZFF_Y2[2:2]),.I4(ZFF_Y2[16:16]),.I5(ZFF_Y2[9:9]),.O(un10_6_axb_8));
defparam desc476.INIT=64'h693CC36996C33C96;
  LUT5 un8_0_8_axb_5_cZ(.I0(ZFF_X2_fast[10:10]),.I1(ZFF_X2_fast[6:6]),.I2(ZFF_X2_fast[0:0]),.I3(ZFF_X2_fast[7:7]),.I4(ZFF_X2_fast[9:9]),.O(un8_0_8_axb_5));
defparam un8_0_8_axb_5_cZ.INIT=32'hA596965A;
  LUT2 un7_0_10_o5_16_cZ(.I0(ZFF_X1[6:6]),.I1(ZFF_X1[9:9]),.O(un7_0_10_o5_16));
defparam un7_0_10_o5_16_cZ.INIT=4'hB;
  LUT6 un8_0_0_axb_20_cZ(.I0(un8_0_8[19:19]),.I1(un8_0_8[20:20]),.I2(un8_0_9[19:19]),.I3(un8_0_9[20:20]),.I4(un8_0_6[19:19]),.I5(un8_0_6[20:20]),.O(un8_0_0_axb_20));
defparam un8_0_0_axb_20_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un6_0_0_axb_16_cZ(.I0(un6_0_9[15:15]),.I1(un6_0_8[15:15]),.I2(un6_0_8[16:16]),.I3(un6_0_9[16:16]),.I4(un6_0_6[15:15]),.I5(un6_0_6[16:16]),.O(un6_0_0_axb_16));
defparam un6_0_0_axb_16_cZ.INIT=64'h1EE17887E11E8778;
  LUT5 un10_axb_21_cZ(.I0(ZFF_Y2[17:17]),.I1(un10_8[26:26]),.I2(un10_8[27:27]),.I3(un10_6[26:26]),.I4(un10_6[27:27]),.O(un10_axb_21));
defparam un10_axb_21_cZ.INIT=32'h871E78E1;
  LUT6 un9_6_78_RNITVCD1(.I0(un9_11_fast[26:26]),.I1(un9_11_22_rep1),.I2(ZFF_Y1_5_rep1),.I3(ZFF_Y1_16_rep1),.I4(ZFF_Y1_4_rep1),.I5(un9_6_78),.O(un9_6_0_axb_22));
defparam un9_6_78_RNITVCD1.INIT=64'h6969699669969696;
  LUT6 un7_0_0_axb_19_cZ(.I0(un7_0_10[18:18]),.I1(un7_0_6[18:18]),.I2(un7_0_6[19:19]),.I3(un7_0_10[19:19]),.I4(un7_0_8[18:18]),.I5(un7_0_8[19:19]),.O(un7_0_0_axb_19));
defparam un7_0_0_axb_19_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 un9_axb_11_cZ(.I0(un9_10[12:12]),.I1(un9_8[12:12]),.I2(un9_8[13:13]),.I3(un9_10[13:13]),.I4(un9_6[12:12]),.I5(un9_6[13:13]),.O(un9_axb_11));
defparam un9_axb_11_cZ.INIT=64'h1EE17887E11E8778;
  LUT6 un8_0_0_axb_16_cZ(.I0(un8_0_9[15:15]),.I1(un8_0_8[15:15]),.I2(un8_0_8[16:16]),.I3(un8_0_9[16:16]),.I4(un8_0_6[15:15]),.I5(un8_0_6[16:16]),.O(un8_0_0_axb_16));
defparam un8_0_0_axb_16_cZ.INIT=64'h1EE17887E11E8778;
  LUT5 un10_axb_20_cZ(.I0(ZFF_Y2[17:17]),.I1(un10_8[25:25]),.I2(un10_8[26:26]),.I3(un10_6[25:25]),.I4(un10_6[26:26]),.O(un10_axb_20));
defparam un10_axb_20_cZ.INIT=32'h871E78E1;
  LUT5 un10_axb_22_cZ(.I0(ZFF_Y2[17:17]),.I1(un10_8[27:27]),.I2(un10_8[28:28]),.I3(un10_6[27:27]),.I4(un10_6[28:28]),.O(un10_axb_22));
defparam un10_axb_22_cZ.INIT=32'h871E78E1;
  LUT6 un9_axb_37_cZ(.I0(un9_8[39:39]),.I1(un9_10[38:38]),.I2(un9_10[39:39]),.I3(un9_8[38:38]),.I4(un9_6[38:38]),.I5(un9_6[39:39]),.O(un9_axb_37));
defparam un9_axb_37_cZ.INIT=64'h5A6969A5A596965A;
  MUXCY_L un9_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un9_ac0_105),.LO(un9_cry_0_cy));
  MUXCY_L un10_8_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un10_8_ac0_5),.LO(un10_8_cry_0_cy));
  LUT5 un9_6_0_cry_5_RNO_0_cZ(.I0(un9_10_fast[8:8]),.I1(ZFF_Y1_fast[3:3]),.I2(ZFF_Y1_fast[4:4]),.I3(un9_8_fast[7:7]),.I4(ZFF_Y1_fast[5:5]),.O(un9_6_0_cry_5_RNO_0));
defparam un9_6_0_cry_5_RNO_0_cZ.INIT=32'hAAAB5554;
  LUT5 un10_6_cry_0_RNO_0_cZ(.I0(ZFF_Y2_fast[8:8]),.I1(ZFF_Y2[0:0]),.I2(ZFF_Y2[2:2]),.I3(ZFF_Y2[1:1]),.I4(ZFF_Y2[9:9]),.O(un10_6_cry_0_RNO_0));
defparam un10_6_cry_0_RNO_0_cZ.INIT=32'hD42B2BD4;
  LUT2 un8_0_0_o5_12_cZ(.I0(un8_0_8[12:12]),.I1(un8_0_6[12:12]),.O(un8_0_0_o5_12));
defparam un8_0_0_o5_12_cZ.INIT=4'h8;
  LUT2 un8_0_0_o5_13_cZ(.I0(un8_0_8[13:13]),.I1(un8_0_6[13:13]),.O(un8_0_0_o5_13));
defparam un8_0_0_o5_13_cZ.INIT=4'h8;
  LUT2 un8_0_0_o5_14_cZ(.I0(un8_0_8[14:14]),.I1(un8_0_6[14:14]),.O(un8_0_0_o5_14));
defparam un8_0_0_o5_14_cZ.INIT=4'h8;
  LUT2_L un9_6_78_cZ(.I0(ZFF_Y1_fast[15:15]),.I1(ZFF_Y1_3_rep1),.LO(un9_6_78));
defparam un9_6_78_cZ.INIT=4'h8;
  LUT2 un6_0_0_o5_12_cZ(.I0(un6_0_8[12:12]),.I1(un6_0_6[12:12]),.O(un6_0_0_o5_12));
defparam un6_0_0_o5_12_cZ.INIT=4'h8;
  LUT2 un6_0_0_o5_13_cZ(.I0(un6_0_8[13:13]),.I1(un6_0_6[13:13]),.O(un6_0_0_o5_13));
defparam un6_0_0_o5_13_cZ.INIT=4'h8;
  LUT2 un6_0_0_o5_14_cZ(.I0(un6_0_8[14:14]),.I1(un6_0_6[14:14]),.O(un6_0_0_o5_14));
defparam un6_0_0_o5_14_cZ.INIT=4'h8;
  LUT2 Y_out_double_2_4_axb_17_cZ(.I0(pgZFF_X2[16:16]),.I1(Y_out_double_2_7[17:17]),.O(Y_out_double_2_4_axb_17));
defparam Y_out_double_2_4_axb_17_cZ.INIT=4'h6;
  LUT2_L un9_11_axb_6(.I0(un9_10_8_rep1),.I1(ZFF_Y1_15_rep1),.LO(un9_11[27:27]));
defparam un9_11_axb_6.INIT=4'h6;
  LUT2 un8_0_9_axb_0(.I0(ZFF_X2_fast[8:8]),.I1(ZFF_X2_fast[7:7]),.O(un8_0_9[15:15]));
defparam un8_0_9_axb_0.INIT=4'h6;
  LUT2 un6_0_9_axb_0(.I0(ZFF_X0_fast[7:7]),.I1(ZFF_X0_fast[8:8]),.O(un6_0_9[15:15]));
defparam un6_0_9_axb_0.INIT=4'h6;
  LUT1 Y_out_double_2_7_axb_16_cZ(.I0(pgZFF_X0[16:16]),.O(Y_out_double_2_7_axb_16));
defparam Y_out_double_2_7_axb_16_cZ.INIT=2'h2;
  LUT2_L Y_out_double_2_axb_17_cZ(.I0(Y_out_double_2_6[17:17]),.I1(Y_out_double_2_4[17:17]),.LO(Y_out_double_2_axb_17));
defparam Y_out_double_2_axb_17_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_16_cZ(.I0(Y_out_double_2_6[16:16]),.I1(Y_out_double_2_4[16:16]),.LO(Y_out_double_2_axb_16));
defparam Y_out_double_2_axb_16_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_15_cZ(.I0(Y_out_double_2_6[15:15]),.I1(Y_out_double_2_4[15:15]),.LO(Y_out_double_2_axb_15));
defparam Y_out_double_2_axb_15_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_14_cZ(.I0(Y_out_double_2_6[14:14]),.I1(Y_out_double_2_4[14:14]),.LO(Y_out_double_2_axb_14));
defparam Y_out_double_2_axb_14_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_13_cZ(.I0(Y_out_double_2_6[13:13]),.I1(Y_out_double_2_4[13:13]),.LO(Y_out_double_2_axb_13));
defparam Y_out_double_2_axb_13_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_12_cZ(.I0(Y_out_double_2_6[12:12]),.I1(Y_out_double_2_4[12:12]),.LO(Y_out_double_2_axb_12));
defparam Y_out_double_2_axb_12_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_11_cZ(.I0(Y_out_double_2_6[11:11]),.I1(Y_out_double_2_4[11:11]),.LO(Y_out_double_2_axb_11));
defparam Y_out_double_2_axb_11_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_10_cZ(.I0(Y_out_double_2_6[10:10]),.I1(Y_out_double_2_4[10:10]),.LO(Y_out_double_2_axb_10));
defparam Y_out_double_2_axb_10_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_9_cZ(.I0(Y_out_double_2_6[9:9]),.I1(Y_out_double_2_4[9:9]),.LO(Y_out_double_2_axb_9));
defparam Y_out_double_2_axb_9_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_8_cZ(.I0(Y_out_double_2_6[8:8]),.I1(Y_out_double_2_4[8:8]),.LO(Y_out_double_2_axb_8));
defparam Y_out_double_2_axb_8_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_7_cZ(.I0(Y_out_double_2_6[7:7]),.I1(Y_out_double_2_4[7:7]),.LO(Y_out_double_2_axb_7));
defparam Y_out_double_2_axb_7_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_6_cZ(.I0(Y_out_double_2_6[6:6]),.I1(Y_out_double_2_4[6:6]),.LO(Y_out_double_2_axb_6));
defparam Y_out_double_2_axb_6_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_5_cZ(.I0(Y_out_double_2_6[5:5]),.I1(Y_out_double_2_4[5:5]),.LO(Y_out_double_2_axb_5));
defparam Y_out_double_2_axb_5_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_4_cZ(.I0(Y_out_double_2_6[4:4]),.I1(Y_out_double_2_4[4:4]),.LO(Y_out_double_2_axb_4));
defparam Y_out_double_2_axb_4_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_3_cZ(.I0(Y_out_double_2_6[3:3]),.I1(Y_out_double_2_4[3:3]),.LO(Y_out_double_2_axb_3));
defparam Y_out_double_2_axb_3_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_2_cZ(.I0(Y_out_double_2_6[2:2]),.I1(Y_out_double_2_4[2:2]),.LO(Y_out_double_2_axb_2));
defparam Y_out_double_2_axb_2_cZ.INIT=4'h6;
  LUT2_L Y_out_double_2_axb_1_cZ(.I0(Y_out_double_2_6[1:1]),.I1(Y_out_double_2_4[1:1]),.LO(Y_out_double_2_axb_1));
defparam Y_out_double_2_axb_1_cZ.INIT=4'h6;
  LUT1 un10_8_axb_28_cZ(.I0(ZFF_Y2[17:17]),.O(un10_8_axb_28));
defparam un10_8_axb_28_cZ.INIT=2'h2;
  LUT2 un7_0_0_axb_45_cZ(.I0(ZFF_X1[16:16]),.I1(un7_0_10[45:45]),.O(un7_0_0_axb_45));
defparam un7_0_0_axb_45_cZ.INIT=4'h6;
  LUT1 desc477(.I0(un10_8[47:47]),.O(un10_8_i[47:47]));
defparam desc477.INIT=2'h1;
  LUT2 un9_10_axb_0(.I0(un9_10_fast[8:8]),.I1(un9_8_7_rep1),.O(un9_10[12:12]));
defparam un9_10_axb_0.INIT=4'h6;
  LUT2 un8_0_8_o5_11_cZ(.I0(ZFF_X2[6:6]),.I1(ZFF_X2[1:1]),.O(un8_0_8_o5_11));
defparam un8_0_8_o5_11_cZ.INIT=4'hD;
  LUT2 un6_0_8_o5_11_cZ(.I0(ZFF_X0[1:1]),.I1(ZFF_X0[6:6]),.O(un6_0_8_o5_11));
defparam un6_0_8_o5_11_cZ.INIT=4'hB;
  LUT2 un7_0_6_o5_16_cZ(.I0(ZFF_X1[2:2]),.I1(ZFF_X1[9:9]),.O(un7_0_6_o5_16));
defparam un7_0_6_o5_16_cZ.INIT=4'hD;
  LUT2 un7_0_6_o5_17_cZ(.I0(ZFF_X1[3:3]),.I1(ZFF_X1[10:10]),.O(un7_0_6_o5_17));
defparam un7_0_6_o5_17_cZ.INIT=4'hD;
  LUT2 un7_0_6_o5_18_cZ(.I0(ZFF_X1[4:4]),.I1(ZFF_X1[11:11]),.O(un7_0_6_o5_18));
defparam un7_0_6_o5_18_cZ.INIT=4'hD;
  LUT2 un7_0_6_o5_19_cZ(.I0(ZFF_X1[5:5]),.I1(ZFF_X1[12:12]),.O(un7_0_6_o5_19));
defparam un7_0_6_o5_19_cZ.INIT=4'hD;
  LUT2 un10_o5_23_cZ(.I0(un10_8[29:29]),.I1(un10_6[29:29]),.O(un10_o5_23));
defparam un10_o5_23_cZ.INIT=4'hE;
  LUT2 un10_o5_24_cZ(.I0(un10_8[30:30]),.I1(un10_6[30:30]),.O(un10_o5_24));
defparam un10_o5_24_cZ.INIT=4'hE;
  LUT2 un10_o5_25_cZ(.I0(un10_8[31:31]),.I1(un10_6[31:31]),.O(un10_o5_25));
defparam un10_o5_25_cZ.INIT=4'hE;
  LUT2 un10_o5_26_cZ(.I0(un10_8[32:32]),.I1(un10_6[32:32]),.O(un10_o5_26));
defparam un10_o5_26_cZ.INIT=4'hE;
  LUT2 un10_o5_27_cZ(.I0(un10_8[33:33]),.I1(un10_6[33:33]),.O(un10_o5_27));
defparam un10_o5_27_cZ.INIT=4'hE;
  LUT2 un9_8_o5_14_cZ(.I0(un9_8[6:6]),.I1(ZFF_Y1[8:8]),.O(un9_8_o5_14));
defparam un9_8_o5_14_cZ.INIT=4'hB;
  LUT2 un9_8_o5_15_cZ(.I0(ZFF_Y1[9:9]),.I1(un9_8[7:7]),.O(un9_8_o5_15));
defparam un9_8_o5_15_cZ.INIT=4'hD;
  LUT2 un7_0_10_o5_15_cZ(.I0(ZFF_X1[5:5]),.I1(ZFF_X1[8:8]),.O(un7_0_10_o5_15));
defparam un7_0_10_o5_15_cZ.INIT=4'hB;
  LUT2 un7_0_10_o5_17_cZ(.I0(ZFF_X1[10:10]),.I1(ZFF_X1[7:7]),.O(un7_0_10_o5_17));
defparam un7_0_10_o5_17_cZ.INIT=4'hD;
  LUT2 un7_0_10_o5_18_cZ(.I0(ZFF_X1[8:8]),.I1(ZFF_X1[11:11]),.O(un7_0_10_o5_18));
defparam un7_0_10_o5_18_cZ.INIT=4'hB;
  LUT2 desc478(.I0(ZFF_X1[8:8]),.I1(ZFF_X1[11:11]),.O(un7_0_10_i_i[17:17]));
defparam desc478.INIT=4'h9;
  LUT3 un9_axb_45_cZ(.I0(un9_8[46:46]),.I1(un9_6[47:47]),.I2(un9_6[46:46]),.O(un9_axb_45));
defparam un9_axb_45_cZ.INIT=8'h93;
  LUT2 un8_0_0_axb_43_cZ(.I0(ZFF_X2[16:16]),.I1(un8_0_9[42:42]),.O(un8_0_0_axb_43));
defparam un8_0_0_axb_43_cZ.INIT=4'hB;
  LUT2 un6_0_0_axb_43_cZ(.I0(ZFF_X0[16:16]),.I1(un6_0_9[42:42]),.O(un6_0_0_axb_43));
defparam un6_0_0_axb_43_cZ.INIT=4'hB;
  LUT3 un7_0_10_o5_14_cZ(.I0(ZFF_X1_fast[16:16]),.I1(ZFF_X1[4:4]),.I2(ZFF_X1[7:7]),.O(un7_0_10_o5_14));
defparam un7_0_10_o5_14_cZ.INIT=8'h8E;
  LUT3 un6_0_0_o5_37_cZ(.I0(ZFF_X0[16:16]),.I1(un6_0_8[37:37]),.I2(un6_0_9[37:37]),.O(un6_0_0_o5_37));
defparam un6_0_0_o5_37_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_27_cZ(.I0(un6_0_8[27:27]),.I1(un6_0_9[27:27]),.I2(un6_0_6[27:27]),.O(un6_0_0_o5_27));
defparam un6_0_0_o5_27_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_26_cZ(.I0(un6_0_8[26:26]),.I1(un6_0_9[26:26]),.I2(un6_0_6[26:26]),.O(un6_0_0_o5_26));
defparam un6_0_0_o5_26_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_25_cZ(.I0(un6_0_8[25:25]),.I1(un6_0_9[25:25]),.I2(un6_0_6[25:25]),.O(un6_0_0_o5_25));
defparam un6_0_0_o5_25_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_24_cZ(.I0(un6_0_8[24:24]),.I1(un6_0_9[24:24]),.I2(un6_0_6[24:24]),.O(un6_0_0_o5_24));
defparam un6_0_0_o5_24_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_23_cZ(.I0(un6_0_8[23:23]),.I1(un6_0_9[23:23]),.I2(un6_0_6[23:23]),.O(un6_0_0_o5_23));
defparam un6_0_0_o5_23_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_22_cZ(.I0(un6_0_8[22:22]),.I1(un6_0_9[22:22]),.I2(un6_0_6[22:22]),.O(un6_0_0_o5_22));
defparam un6_0_0_o5_22_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_21_cZ(.I0(un6_0_8[21:21]),.I1(un6_0_9[21:21]),.I2(un6_0_6[21:21]),.O(un6_0_0_o5_21));
defparam un6_0_0_o5_21_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_20_cZ(.I0(un6_0_8[20:20]),.I1(un6_0_9[20:20]),.I2(un6_0_6[20:20]),.O(un6_0_0_o5_20));
defparam un6_0_0_o5_20_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_19_cZ(.I0(un6_0_8[19:19]),.I1(un6_0_9[19:19]),.I2(un6_0_6[19:19]),.O(un6_0_0_o5_19));
defparam un6_0_0_o5_19_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_18_cZ(.I0(un6_0_8[18:18]),.I1(un6_0_9[18:18]),.I2(un6_0_6[18:18]),.O(un6_0_0_o5_18));
defparam un6_0_0_o5_18_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_17_cZ(.I0(un6_0_8[17:17]),.I1(un6_0_9[17:17]),.I2(un6_0_6[17:17]),.O(un6_0_0_o5_17));
defparam un6_0_0_o5_17_cZ.INIT=8'hE8;
  LUT3 un6_0_0_o5_16_cZ(.I0(un6_0_8[16:16]),.I1(un6_0_9[16:16]),.I2(un6_0_6[16:16]),.O(un6_0_0_o5_16));
defparam un6_0_0_o5_16_cZ.INIT=8'hE8;
  LUT3 un9_o5_39_cZ(.I0(un9_8[41:41]),.I1(un9_10[41:41]),.I2(un9_6[41:41]),.O(un9_o5_39));
defparam un9_o5_39_cZ.INIT=8'hE8;
  LUT3 un9_o5_38_cZ(.I0(un9_8[40:40]),.I1(un9_10[40:40]),.I2(un9_6[40:40]),.O(un9_o5_38));
defparam un9_o5_38_cZ.INIT=8'hE8;
  LUT3 un9_o5_37_cZ(.I0(un9_8[39:39]),.I1(un9_10[39:39]),.I2(un9_6[39:39]),.O(un9_o5_37));
defparam un9_o5_37_cZ.INIT=8'hE8;
  LUT3 un9_o5_35_cZ(.I0(un9_8[37:37]),.I1(un9_10[37:37]),.I2(un9_6[37:37]),.O(un9_o5_35));
defparam un9_o5_35_cZ.INIT=8'hE8;
  LUT3 un9_o5_34_cZ(.I0(un9_8[36:36]),.I1(un9_10[36:36]),.I2(un9_6[36:36]),.O(un9_o5_34));
defparam un9_o5_34_cZ.INIT=8'hE8;
  LUT3 un9_o5_33_cZ(.I0(un9_8[35:35]),.I1(un9_10[35:35]),.I2(un9_6[35:35]),.O(un9_o5_33));
defparam un9_o5_33_cZ.INIT=8'hE8;
  LUT3 un9_o5_32_cZ(.I0(un9_8[34:34]),.I1(un9_10[34:34]),.I2(un9_6[34:34]),.O(un9_o5_32));
defparam un9_o5_32_cZ.INIT=8'hE8;
  LUT3 un9_o5_31_cZ(.I0(un9_8[33:33]),.I1(un9_10[33:33]),.I2(un9_6[33:33]),.O(un9_o5_31));
defparam un9_o5_31_cZ.INIT=8'hE8;
  LUT3 un9_o5_30_cZ(.I0(un9_8[32:32]),.I1(un9_10[32:32]),.I2(un9_6[32:32]),.O(un9_o5_30));
defparam un9_o5_30_cZ.INIT=8'hE8;
  LUT3 un9_o5_29_cZ(.I0(un9_8[31:31]),.I1(un9_10[31:31]),.I2(un9_6[31:31]),.O(un9_o5_29));
defparam un9_o5_29_cZ.INIT=8'hE8;
  LUT3 un9_o5_28_cZ(.I0(un9_8[30:30]),.I1(un9_10[30:30]),.I2(un9_6[30:30]),.O(un9_o5_28));
defparam un9_o5_28_cZ.INIT=8'hE8;
  LUT3 un9_o5_27_cZ(.I0(un9_8[29:29]),.I1(un9_10[29:29]),.I2(un9_6[29:29]),.O(un9_o5_27));
defparam un9_o5_27_cZ.INIT=8'hE8;
  LUT3 un9_o5_26_cZ(.I0(un9_8[28:28]),.I1(un9_10[28:28]),.I2(un9_6[28:28]),.O(un9_o5_26));
defparam un9_o5_26_cZ.INIT=8'hE8;
  LUT3 un9_o5_25_cZ(.I0(un9_8[27:27]),.I1(un9_10[27:27]),.I2(un9_6[27:27]),.O(un9_o5_25));
defparam un9_o5_25_cZ.INIT=8'hE8;
  LUT3 un9_o5_24_cZ(.I0(un9_8[26:26]),.I1(un9_10[26:26]),.I2(un9_6[26:26]),.O(un9_o5_24));
defparam un9_o5_24_cZ.INIT=8'hE8;
  LUT3 un9_o5_23_cZ(.I0(un9_8[25:25]),.I1(un9_10[25:25]),.I2(un9_6[25:25]),.O(un9_o5_23));
defparam un9_o5_23_cZ.INIT=8'hE8;
  LUT3 un9_o5_22_cZ(.I0(un9_8[24:24]),.I1(un9_10[24:24]),.I2(un9_6[24:24]),.O(un9_o5_22));
defparam un9_o5_22_cZ.INIT=8'hE8;
  LUT3 un9_o5_21_cZ(.I0(un9_8[23:23]),.I1(un9_10[23:23]),.I2(un9_6[23:23]),.O(un9_o5_21));
defparam un9_o5_21_cZ.INIT=8'hE8;
  LUT3 un9_o5_20_cZ(.I0(un9_8[22:22]),.I1(un9_10[22:22]),.I2(un9_6[22:22]),.O(un9_o5_20));
defparam un9_o5_20_cZ.INIT=8'hE8;
  LUT3 un9_o5_19_cZ(.I0(un9_8[21:21]),.I1(un9_10[21:21]),.I2(un9_6[21:21]),.O(un9_o5_19));
defparam un9_o5_19_cZ.INIT=8'hE8;
  LUT3 un9_o5_18_cZ(.I0(un9_8[20:20]),.I1(un9_10[20:20]),.I2(un9_6[20:20]),.O(un9_o5_18));
defparam un9_o5_18_cZ.INIT=8'hE8;
  LUT3 un9_o5_17_cZ(.I0(un9_8[19:19]),.I1(un9_10[19:19]),.I2(un9_6[19:19]),.O(un9_o5_17));
defparam un9_o5_17_cZ.INIT=8'hE8;
  LUT3 un9_o5_16_cZ(.I0(un9_8[18:18]),.I1(un9_10[18:18]),.I2(un9_6[18:18]),.O(un9_o5_16));
defparam un9_o5_16_cZ.INIT=8'hE8;
  LUT3 un9_o5_15_cZ(.I0(un9_8[17:17]),.I1(un9_10[17:17]),.I2(un9_6[17:17]),.O(un9_o5_15));
defparam un9_o5_15_cZ.INIT=8'hE8;
  LUT3 un9_o5_14_cZ(.I0(un9_8[16:16]),.I1(un9_10[16:16]),.I2(un9_6[16:16]),.O(un9_o5_14));
defparam un9_o5_14_cZ.INIT=8'hE8;
  LUT3 un9_o5_13_cZ(.I0(un9_8[15:15]),.I1(un9_10[15:15]),.I2(un9_6[15:15]),.O(un9_o5_13));
defparam un9_o5_13_cZ.INIT=8'hE8;
  LUT3 un9_o5_12_cZ(.I0(un9_8[14:14]),.I1(un9_10[14:14]),.I2(un9_6[14:14]),.O(un9_o5_12));
defparam un9_o5_12_cZ.INIT=8'hE8;
  LUT3 un9_o5_11_cZ(.I0(un9_8[13:13]),.I1(un9_10[13:13]),.I2(un9_6[13:13]),.O(un9_o5_11));
defparam un9_o5_11_cZ.INIT=8'hE8;
  LUT3 un9_o5_9_cZ(.I0(ZFF_Y1[6:6]),.I1(un9_8[11:11]),.I2(un9_6[11:11]),.O(un9_o5_9));
defparam un9_o5_9_cZ.INIT=8'hE8;
  LUT3 un9_o5_8_cZ(.I0(ZFF_Y1[5:5]),.I1(un9_8[10:10]),.I2(un9_6[10:10]),.O(un9_o5_8));
defparam un9_o5_8_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_37_cZ(.I0(ZFF_X2[16:16]),.I1(un8_0_8[37:37]),.I2(un8_0_9[37:37]),.O(un8_0_0_o5_37));
defparam un8_0_0_o5_37_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_27_cZ(.I0(un8_0_8[27:27]),.I1(un8_0_9[27:27]),.I2(un8_0_6[27:27]),.O(un8_0_0_o5_27));
defparam un8_0_0_o5_27_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_26_cZ(.I0(un8_0_8[26:26]),.I1(un8_0_9[26:26]),.I2(un8_0_6[26:26]),.O(un8_0_0_o5_26));
defparam un8_0_0_o5_26_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_25_cZ(.I0(un8_0_8[25:25]),.I1(un8_0_9[25:25]),.I2(un8_0_6[25:25]),.O(un8_0_0_o5_25));
defparam un8_0_0_o5_25_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_24_cZ(.I0(un8_0_8[24:24]),.I1(un8_0_9[24:24]),.I2(un8_0_6[24:24]),.O(un8_0_0_o5_24));
defparam un8_0_0_o5_24_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_23_cZ(.I0(un8_0_8[23:23]),.I1(un8_0_9[23:23]),.I2(un8_0_6[23:23]),.O(un8_0_0_o5_23));
defparam un8_0_0_o5_23_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_22_cZ(.I0(un8_0_8[22:22]),.I1(un8_0_9[22:22]),.I2(un8_0_6[22:22]),.O(un8_0_0_o5_22));
defparam un8_0_0_o5_22_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_21_cZ(.I0(un8_0_8[21:21]),.I1(un8_0_9[21:21]),.I2(un8_0_6[21:21]),.O(un8_0_0_o5_21));
defparam un8_0_0_o5_21_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_20_cZ(.I0(un8_0_8[20:20]),.I1(un8_0_9[20:20]),.I2(un8_0_6[20:20]),.O(un8_0_0_o5_20));
defparam un8_0_0_o5_20_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_19_cZ(.I0(un8_0_8[19:19]),.I1(un8_0_9[19:19]),.I2(un8_0_6[19:19]),.O(un8_0_0_o5_19));
defparam un8_0_0_o5_19_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_18_cZ(.I0(un8_0_8[18:18]),.I1(un8_0_9[18:18]),.I2(un8_0_6[18:18]),.O(un8_0_0_o5_18));
defparam un8_0_0_o5_18_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_17_cZ(.I0(un8_0_8[17:17]),.I1(un8_0_9[17:17]),.I2(un8_0_6[17:17]),.O(un8_0_0_o5_17));
defparam un8_0_0_o5_17_cZ.INIT=8'hE8;
  LUT3 un8_0_0_o5_16_cZ(.I0(un8_0_8[16:16]),.I1(un8_0_9[16:16]),.I2(un8_0_6[16:16]),.O(un8_0_0_o5_16));
defparam un8_0_0_o5_16_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_32_cZ(.I0(un7_0_6[32:32]),.I1(un7_0_10[32:32]),.I2(un7_0_8[32:32]),.O(un7_0_0_o5_32));
defparam un7_0_0_o5_32_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_31_cZ(.I0(un7_0_6[31:31]),.I1(un7_0_10[31:31]),.I2(un7_0_8[31:31]),.O(un7_0_0_o5_31));
defparam un7_0_0_o5_31_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_30_cZ(.I0(un7_0_6[30:30]),.I1(un7_0_10[30:30]),.I2(un7_0_8[30:30]),.O(un7_0_0_o5_30));
defparam un7_0_0_o5_30_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_29_cZ(.I0(un7_0_6[29:29]),.I1(un7_0_10[29:29]),.I2(un7_0_8[29:29]),.O(un7_0_0_o5_29));
defparam un7_0_0_o5_29_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_28_cZ(.I0(un7_0_6[28:28]),.I1(un7_0_10[28:28]),.I2(un7_0_8[28:28]),.O(un7_0_0_o5_28));
defparam un7_0_0_o5_28_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_27_cZ(.I0(un7_0_6[27:27]),.I1(un7_0_10[27:27]),.I2(un7_0_8[27:27]),.O(un7_0_0_o5_27));
defparam un7_0_0_o5_27_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_26_cZ(.I0(un7_0_6[26:26]),.I1(un7_0_10[26:26]),.I2(un7_0_8[26:26]),.O(un7_0_0_o5_26));
defparam un7_0_0_o5_26_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_25_cZ(.I0(un7_0_6[25:25]),.I1(un7_0_10[25:25]),.I2(un7_0_8[25:25]),.O(un7_0_0_o5_25));
defparam un7_0_0_o5_25_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_24_cZ(.I0(un7_0_6[24:24]),.I1(un7_0_10[24:24]),.I2(un7_0_8[24:24]),.O(un7_0_0_o5_24));
defparam un7_0_0_o5_24_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_23_cZ(.I0(un7_0_6[23:23]),.I1(un7_0_10[23:23]),.I2(un7_0_8[23:23]),.O(un7_0_0_o5_23));
defparam un7_0_0_o5_23_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_22_cZ(.I0(un7_0_6[22:22]),.I1(un7_0_10[22:22]),.I2(un7_0_8[22:22]),.O(un7_0_0_o5_22));
defparam un7_0_0_o5_22_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_21_cZ(.I0(un7_0_6[21:21]),.I1(un7_0_10[21:21]),.I2(un7_0_8[21:21]),.O(un7_0_0_o5_21));
defparam un7_0_0_o5_21_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_20_cZ(.I0(un7_0_6[20:20]),.I1(un7_0_10[20:20]),.I2(un7_0_8[20:20]),.O(un7_0_0_o5_20));
defparam un7_0_0_o5_20_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_19_cZ(.I0(un7_0_6[19:19]),.I1(un7_0_10[19:19]),.I2(un7_0_8[19:19]),.O(un7_0_0_o5_19));
defparam un7_0_0_o5_19_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_16_cZ(.I0(ZFF_X1[13:13]),.I1(un7_0_6[16:16]),.I2(un7_0_8[16:16]),.O(un7_0_0_o5_16));
defparam un7_0_0_o5_16_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_15_cZ(.I0(ZFF_X1[12:12]),.I1(un7_0_6[15:15]),.I2(un7_0_8[15:15]),.O(un7_0_0_o5_15));
defparam un7_0_0_o5_15_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_14_cZ(.I0(ZFF_X1[11:11]),.I1(un7_0_6[14:14]),.I2(un7_0_8[14:14]),.O(un7_0_0_o5_14));
defparam un7_0_0_o5_14_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_13_cZ(.I0(ZFF_X1[7:7]),.I1(un7_0_6[13:13]),.I2(un7_0_8[13:13]),.O(un7_0_0_o5_13));
defparam un7_0_0_o5_13_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_12_cZ(.I0(ZFF_X1[6:6]),.I1(un7_0_6[12:12]),.I2(un7_0_8[12:12]),.O(un7_0_0_o5_12));
defparam un7_0_0_o5_12_cZ.INIT=8'hE8;
  LUT3 un7_0_0_o5_11_cZ(.I0(ZFF_X1[2:2]),.I1(un7_0_6[11:11]),.I2(un7_0_8[11:11]),.O(un7_0_0_o5_11));
defparam un7_0_0_o5_11_cZ.INIT=8'hE8;
  LUT3 un7_0_6_o5_15_cZ(.I0(ZFF_X1_1_rep1),.I1(ZFF_X1_8_rep1),.I2(ZFF_X1_fast[16:16]),.O(un7_0_6_o5_15));
defparam un7_0_6_o5_15_cZ.INIT=8'h4D;
  LUT3 un6_0_8_o5_4_cZ(.I0(ZFF_X0_7_rep1),.I1(ZFF_X0_fast[6:6]),.I2(ZFF_X0_fast[9:9]),.O(un6_0_8_o5_4));
defparam un6_0_8_o5_4_cZ.INIT=8'hE8;
  LUT3 un8_0_8_o5_4_cZ(.I0(ZFF_X2_fast[6:6]),.I1(ZFF_X2_fast[7:7]),.I2(ZFF_X2_fast[9:9]),.O(un8_0_8_o5_4));
defparam un8_0_8_o5_4_cZ.INIT=8'hE8;
  LUT4 desc479(.I0(sample_trig),.I1(q_reg_i_1[1:1]),.I2(q_reg_i_1[2:2]),.I3(state_reg),.O(state_next));
defparam desc479.INIT=16'hFCAA;
  LUT5 un10_axb_4_cZ(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[3:3]),.I3(ZFF_Y2[1:1]),.I4(un10_6[10:10]),.O(un10_axb_4));
defparam un10_axb_4_cZ.INIT=32'hCCC63339;
  LUT6 desc480(.I0(q_reg[2:2]),.I1(q_reg[1:1]),.I2(q_reg[0:0]),.I3(q_reg_i_1[1:1]),.I4(q_reg_i_1[2:2]),.I5(state_reg),.O(q_next[2:2]));
defparam desc480.INIT=64'h6A6A6A00AAAAAAAA;
  LUT6_L state_reg_ret_RNO(.I0(q_reg[2:2]),.I1(q_reg[1:1]),.I2(q_reg[0:0]),.I3(q_reg_i_1[1:1]),.I4(q_reg_i_1[2:2]),.I5(state_reg),.LO(q_next_i[2:2]));
defparam state_reg_ret_RNO.INIT=64'h959595FF55555555;
  LUT5 un8_0_0_axb_39_cZ(.I0(ZFF_X2[16:16]),.I1(un8_0_8[39:39]),.I2(un8_0_9[38:38]),.I3(un8_0_9[39:39]),.I4(un8_0_8[38:38]),.O(un8_0_0_axb_39));
defparam un8_0_0_axb_39_cZ.INIT=32'h936CC936;
  LUT5 un6_0_0_axb_39_cZ(.I0(ZFF_X0[16:16]),.I1(un6_0_8[39:39]),.I2(un6_0_9[38:38]),.I3(un6_0_9[39:39]),.I4(un6_0_8[38:38]),.O(un6_0_0_axb_39));
defparam un6_0_0_axb_39_cZ.INIT=32'h936CC936;
  LUT5 un8_0_9_s_25_RNIE09P1(.I0(ZFF_X2[16:16]),.I1(un8_0_9[38:38]),.I2(un8_0_9[39:39]),.I3(un8_0_9[40:40]),.I4(un8_0_8[38:38]),.O(N_1128_i));
defparam un8_0_9_s_25_RNIE09P1.INIT=32'h807FE01F;
  LUT5 un6_0_9_s_25_RNI4CK41(.I0(ZFF_X0[16:16]),.I1(un6_0_9[38:38]),.I2(un6_0_9[39:39]),.I3(un6_0_9[40:40]),.I4(un6_0_8[38:38]),.O(N_2007_i));
defparam un6_0_9_s_25_RNI4CK41.INIT=32'h807FE01F;
  LUT6 un8_0_0_o5_41_cZ(.I0(ZFF_X2[16:16]),.I1(un8_0_9[41:41]),.I2(un8_0_9[38:38]),.I3(un8_0_9[39:39]),.I4(un8_0_9[40:40]),.I5(un8_0_8[38:38]),.O(un8_0_0_o5_41));
defparam un8_0_0_o5_41_cZ.INIT=64'hECCCCCCCFECCCCCC;
  LUT6 un6_0_0_o5_41_cZ(.I0(ZFF_X0[16:16]),.I1(un6_0_9[41:41]),.I2(un6_0_9[38:38]),.I3(un6_0_9[39:39]),.I4(un6_0_9[40:40]),.I5(un6_0_8[38:38]),.O(un6_0_0_o5_41));
defparam un6_0_0_o5_41_cZ.INIT=64'hECCCCCCCFECCCCCC;
  LUT6_L un7_q_reg_0_ac0_3(.I0(q_reg[2:2]),.I1(q_reg[1:1]),.I2(q_reg[0:0]),.I3(q_reg_i_1[1:1]),.I4(q_reg_i_1[2:2]),.I5(state_reg),.LO(un7_q_reg_reti));
defparam un7_q_reg_0_ac0_3.INIT=64'h919191FF15151515;
  LUT6 un8_0_0_axb_41_cZ(.I0(ZFF_X2[16:16]),.I1(un8_0_9[41:41]),.I2(un8_0_9[38:38]),.I3(un8_0_9[39:39]),.I4(un8_0_9[40:40]),.I5(un8_0_8[38:38]),.O(un8_0_0_axb_41));
defparam un8_0_0_axb_41_cZ.INIT=64'h93333333C9333333;
  LUT6 un6_0_0_axb_41_cZ(.I0(ZFF_X0[16:16]),.I1(un6_0_9[41:41]),.I2(un6_0_9[38:38]),.I3(un6_0_9[39:39]),.I4(un6_0_9[40:40]),.I5(un6_0_8[38:38]),.O(un6_0_0_axb_41));
defparam un6_0_0_axb_41_cZ.INIT=64'h93333333C9333333;
  LUT4_L state_reg_ret_5_RNO(.I0(state_next),.I1(q_next[0:0]),.I2(q_next[1:1]),.I3(q_next[2:2]),.LO(un1_q_reg_2_reti));
defparam state_reg_ret_5_RNO.INIT=16'h0028;
  LUT4 desc481(.I0(ZFF_X1_fast[15:15]),.I1(ZFF_X1_fast[9:9]),.I2(ZFF_X1_fast[11:11]),.I3(ZFF_X1_fast[8:8]),.O(un7_0_10[18:18]));
defparam desc481.INIT=16'h9996;
  LUT2 un7_0_10_cry_0_RNO_cZ(.I0(ZFF_X1_fast[11:11]),.I1(ZFF_X1_fast[8:8]),.O(un7_0_10_cry_0_RNO));
defparam un7_0_10_cry_0_RNO_cZ.INIT=4'hE;
  LUT2 un7_0_10_cry_1_RNO_cZ(.I0(ZFF_X1_15_rep1),.I1(ZFF_X1[9:9]),.O(un7_0_10_cry_1_RNO));
defparam un7_0_10_cry_1_RNO_cZ.INIT=4'h8;
  LUT2 un7_0_10_cry_12_RNO_cZ(.I0(ZFF_X1[1:1]),.I1(ZFF_X1[16:16]),.O(un7_0_10_cry_12_RNO));
defparam un7_0_10_cry_12_RNO_cZ.INIT=4'h8;
  LUT2 un7_0_10_cry_13_RNO_cZ(.I0(ZFF_X1[2:2]),.I1(ZFF_X1[5:5]),.O(un7_0_10_cry_13_RNO));
defparam un7_0_10_cry_13_RNO_cZ.INIT=4'h2;
  LUT3 un7_0_10_cry_14_RNO_cZ(.I0(ZFF_X1_fast[16:16]),.I1(ZFF_X1[4:4]),.I2(ZFF_X1[7:7]),.O(un7_0_10_cry_14_RNO));
defparam un7_0_10_cry_14_RNO_cZ.INIT=8'h69;
  LUT5 un6_0_9_s_13_RNIJVR91(.I0(un6_0_6[28:28]),.I1(un6_0_8[28:28]),.I2(un6_0_9[28:28]),.I3(un6_0_8[29:29]),.I4(un6_0_9[29:29]),.O(un6_0_0_axb_29));
defparam un6_0_9_s_13_RNIJVR91.INIT=32'hE81717E8;
  LUT2 un6_0_0_cry_29_RNO_cZ(.I0(un6_0_8[29:29]),.I1(un6_0_9[29:29]),.O(un6_0_0_cry_29_RNO));
defparam un6_0_0_cry_29_RNO_cZ.INIT=4'h6;
  LUT2 un6_0_0_cry_30_RNO_cZ(.I0(un6_0_8[29:29]),.I1(un6_0_9[29:29]),.O(un6_0_0_cry_30_RNO));
defparam un6_0_0_cry_30_RNO_cZ.INIT=4'h8;
  LUT2 un6_0_0_cry_31_RNO_cZ(.I0(un6_0_8[30:30]),.I1(un6_0_9[30:30]),.O(un6_0_0_cry_31_RNO));
defparam un6_0_0_cry_31_RNO_cZ.INIT=4'h8;
  LUT2 un6_0_0_cry_32_RNO_cZ(.I0(un6_0_8[31:31]),.I1(un6_0_9[31:31]),.O(un6_0_0_cry_32_RNO));
defparam un6_0_0_cry_32_RNO_cZ.INIT=4'h8;
  LUT2 un6_0_0_cry_33_RNO_cZ(.I0(un6_0_8[32:32]),.I1(un6_0_9[32:32]),.O(un6_0_0_cry_33_RNO));
defparam un6_0_0_cry_33_RNO_cZ.INIT=4'h8;
  LUT2 un6_0_0_cry_34_RNO_cZ(.I0(un6_0_8[33:33]),.I1(un6_0_9[33:33]),.O(un6_0_0_cry_34_RNO));
defparam un6_0_0_cry_34_RNO_cZ.INIT=4'h8;
  LUT2 un6_0_0_cry_35_RNO_cZ(.I0(un6_0_8[34:34]),.I1(un6_0_9[34:34]),.O(un6_0_0_cry_35_RNO));
defparam un6_0_0_cry_35_RNO_cZ.INIT=4'h8;
  LUT2 un6_0_0_cry_36_RNO_cZ(.I0(un6_0_8[35:35]),.I1(un6_0_9[35:35]),.O(un6_0_0_cry_36_RNO));
defparam un6_0_0_cry_36_RNO_cZ.INIT=4'h8;
  LUT5 ZFF_X0_4_rep1_RNIKIE11(.I0(ZFF_X0_2_rep1),.I1(ZFF_X0_4_rep1),.I2(ZFF_X0_3_rep1),.I3(ZFF_X0_1_rep1),.I4(ZFF_X0[9:9]),.O(un6_0_6_axb_4));
defparam ZFF_X0_4_rep1_RNIKIE11.INIT=32'h96666999;
  LUT2 un6_0_6_cry_4_RNO_cZ(.I0(ZFF_X0_3_rep1),.I1(ZFF_X0_1_rep1),.O(un6_0_6_cry_4_RNO));
defparam un6_0_6_cry_4_RNO_cZ.INIT=4'h8;
  LUT3 un6_0_6_cry_5_RNO_cZ(.I0(ZFF_X0[0:0]),.I1(ZFF_X0[10:10]),.I2(ZFF_X0[5:5]),.O(un6_0_6_cry_5_RNO));
defparam un6_0_6_cry_5_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_6_RNO_cZ(.I0(ZFF_X0[1:1]),.I1(ZFF_X0[6:6]),.I2(ZFF_X0[11:11]),.O(un6_0_6_cry_6_RNO));
defparam un6_0_6_cry_6_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_7_RNO_cZ(.I0(ZFF_X0[2:2]),.I1(ZFF_X0[0:0]),.I2(ZFF_X0[12:12]),.O(un6_0_6_cry_7_RNO));
defparam un6_0_6_cry_7_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_8_RNO_cZ(.I0(ZFF_X0[1:1]),.I1(ZFF_X0[3:3]),.I2(ZFF_X0[13:13]),.O(un6_0_6_cry_8_RNO));
defparam un6_0_6_cry_8_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_9_RNO_cZ(.I0(ZFF_X0[4:4]),.I1(ZFF_X0[14:14]),.I2(ZFF_X0[2:2]),.O(un6_0_6_cry_9_RNO));
defparam un6_0_6_cry_9_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_10_RNO_cZ(.I0(ZFF_X0[3:3]),.I1(ZFF_X0[15:15]),.I2(ZFF_X0[5:5]),.O(un6_0_6_cry_10_RNO));
defparam un6_0_6_cry_10_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_11_RNO_cZ(.I0(ZFF_X0[4:4]),.I1(ZFF_X0[6:6]),.I2(ZFF_X0[16:16]),.O(un6_0_6_cry_11_RNO));
defparam un6_0_6_cry_11_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_12_RNO_cZ(.I0(ZFF_X0_16_rep1),.I1(ZFF_X0[7:7]),.I2(ZFF_X0[5:5]),.O(un6_0_6_cry_12_RNO));
defparam un6_0_6_cry_12_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_13_RNO_cZ(.I0(ZFF_X0_16_rep1),.I1(ZFF_X0[6:6]),.I2(ZFF_X0[8:8]),.O(un6_0_6_cry_13_RNO));
defparam un6_0_6_cry_13_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_14_RNO_cZ(.I0(ZFF_X0_16_rep1),.I1(ZFF_X0[7:7]),.I2(ZFF_X0[9:9]),.O(un6_0_6_cry_14_RNO));
defparam un6_0_6_cry_14_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_15_RNO_cZ(.I0(ZFF_X0_16_rep1),.I1(ZFF_X0[10:10]),.I2(ZFF_X0[8:8]),.O(un6_0_6_cry_15_RNO));
defparam un6_0_6_cry_15_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_6_cry_16_RNO_cZ(.I0(ZFF_X0[16:16]),.I1(ZFF_X0[10:10]),.I2(ZFF_X0[8:8]),.O(un6_0_6_cry_16_RNO));
defparam un6_0_6_cry_16_RNO_cZ.INIT=8'hD4;
  LUT3 un6_0_6_cry_17_RNO_cZ(.I0(ZFF_X0[15:15]),.I1(ZFF_X0[10:10]),.I2(ZFF_X0[12:12]),.O(un6_0_6_cry_17_RNO));
defparam un6_0_6_cry_17_RNO_cZ.INIT=8'h96;
  LUT3 un6_0_6_cry_18_RNO_cZ(.I0(ZFF_X0_15_rep1),.I1(ZFF_X0[11:11]),.I2(ZFF_X0[13:13]),.O(un6_0_6_cry_18_RNO));
defparam un6_0_6_cry_18_RNO_cZ.INIT=8'h96;
  LUT5 ZFF_X0_14_rep1_RNI9KV12(.I0(ZFF_X0_14_rep1),.I1(ZFF_X0_15_rep1),.I2(ZFF_X0[12:12]),.I3(ZFF_X0[11:11]),.I4(ZFF_X0[13:13]),.O(un6_0_6_axb_19));
defparam ZFF_X0_14_rep1_RNI9KV12.INIT=32'hA596965A;
  LUT3 un6_0_6_cry_19_RNO_cZ(.I0(ZFF_X0_15_rep1),.I1(ZFF_X0[11:11]),.I2(ZFF_X0[13:13]),.O(un6_0_6_cry_19_RNO));
defparam un6_0_6_cry_19_RNO_cZ.INIT=8'hE8;
  LUT2 un6_0_6_cry_20_RNO_cZ(.I0(ZFF_X0_14_rep1),.I1(ZFF_X0[12:12]),.O(un6_0_6_cry_20_RNO));
defparam un6_0_6_cry_20_RNO_cZ.INIT=4'h8;
  LUT2 un6_0_6_cry_21_RNO(.I0(ZFF_X0[15:15]),.I1(ZFF_X0[13:13]),.O(un6_0_6_43));
defparam un6_0_6_cry_21_RNO.INIT=4'h8;
  LUT5 un9_8_s_34_RNI1A0A1(.I0(un9_10[42:42]),.I1(un9_8[42:42]),.I2(un9_8[43:43]),.I3(un9_6[42:42]),.I4(un9_6[43:43]),.O(un9_axb_41));
defparam un9_8_s_34_RNI1A0A1.INIT=32'hE1871E78;
  LUT2 un9_cry_41_RNO_cZ(.I0(un9_8[43:43]),.I1(un9_6[43:43]),.O(un9_cry_41_RNO));
defparam un9_cry_41_RNO_cZ.INIT=4'h6;
  LUT2 un9_cry_42_RNO_cZ(.I0(un9_8[43:43]),.I1(un9_6[43:43]),.O(un9_cry_42_RNO));
defparam un9_cry_42_RNO_cZ.INIT=4'h8;
  LUT2 un9_cry_43_RNO_cZ(.I0(un9_8[44:44]),.I1(un9_6[44:44]),.O(un9_cry_43_RNO));
defparam un9_cry_43_RNO_cZ.INIT=4'h8;
  LUT2 un9_cry_44_RNO_cZ(.I0(un9_8[45:45]),.I1(un9_6[45:45]),.O(un9_cry_44_RNO));
defparam un9_cry_44_RNO_cZ.INIT=4'h4;
  LUT4 un9_6_0_cry_5_RNO_cZ(.I0(un9_10_fast[8:8]),.I1(ZFF_Y1_fast[3:3]),.I2(ZFF_Y1_fast[4:4]),.I3(un9_8_fast[7:7]),.O(un9_6_0_cry_5_RNO));
defparam un9_6_0_cry_5_RNO_cZ.INIT=16'h0001;
  LUT2 un9_6_0_cry_6_RNO_cZ(.I0(ZFF_Y1_fast[6:6]),.I1(ZFF_Y1_4_rep1),.O(un9_6_0_cry_6_RNO));
defparam un9_6_0_cry_6_RNO_cZ.INIT=4'h6;
  LUT2 un9_6_0_cry_7_RNO_cZ(.I0(ZFF_Y1_fast[7:7]),.I1(ZFF_Y1_5_rep1),.O(un9_6_0_cry_7_RNO));
defparam un9_6_0_cry_7_RNO_cZ.INIT=4'h6;
  LUT2 un9_6_0_cry_8_RNO_cZ(.I0(ZFF_Y1_fast[7:7]),.I1(ZFF_Y1_5_rep1),.O(un9_6_0_cry_8_RNO));
defparam un9_6_0_cry_8_RNO_cZ.INIT=4'h1;
  LUT2 un9_6_0_cry_11_RNO_cZ(.I0(un9_8_6_rep1),.I1(un9_11_fast[23:23]),.O(un9_6_0_cry_11_RNO));
defparam un9_6_0_cry_11_RNO_cZ.INIT=4'h9;
  LUT2 un9_6_0_cry_12_RNO_cZ(.I0(un9_11_24_rep1),.I1(ZFF_Y1_4_rep1),.O(un9_6_0_cry_12_RNO));
defparam un9_6_0_cry_12_RNO_cZ.INIT=4'h9;
  LUT2 un9_6_0_cry_13_RNO_cZ(.I0(ZFF_Y1[5:5]),.I1(un9_11_25_rep1),.O(un9_6_0_cry_13_RNO));
defparam un9_6_0_cry_13_RNO_cZ.INIT=4'h9;
  LUT2 un9_6_0_cry_14_RNO_cZ(.I0(un9_11_26_rep1),.I1(un9_11_24_rep1),.O(un9_6_0_cry_14_RNO));
defparam un9_6_0_cry_14_RNO_cZ.INIT=4'h6;
  LUT2 un9_6_0_cry_15_RNO_cZ(.I0(un9_11_22_rep1),.I1(ZFF_Y1_15_rep1),.O(un9_6_0_cry_15_RNO));
defparam un9_6_0_cry_15_RNO_cZ.INIT=4'h9;
  LUT2 un9_6_0_cry_16_RNO_cZ(.I0(un9_11_23_rep1),.I1(ZFF_Y1_16_rep1),.O(un9_6_0_cry_16_RNO));
defparam un9_6_0_cry_16_RNO_cZ.INIT=4'h9;
  LUT2 un9_6_0_cry_17_RNO_cZ(.I0(ZFF_Y1_17_rep1),.I1(un9_10[8:8]),.O(un9_6_0_cry_17_RNO));
defparam un9_6_0_cry_17_RNO_cZ.INIT=4'h9;
  LUT2 un9_6_0_cry_18_RNO_cZ(.I0(un9_8[6:6]),.I1(ZFF_Y1[17:17]),.O(un9_6_0_cry_18_RNO));
defparam un9_6_0_cry_18_RNO_cZ.INIT=4'h9;
  LUT2 un9_6_0_cry_19_RNO_cZ(.I0(un9_11_23_rep1),.I1(un9_8[7:7]),.O(un9_6_0_cry_19_RNO));
defparam un9_6_0_cry_19_RNO_cZ.INIT=4'h6;
  LUT2 un9_6_0_cry_20_RNO_cZ(.I0(ZFF_Y1_15_rep1),.I1(ZFF_Y1[3:3]),.O(un9_6_0_cry_20_RNO));
defparam un9_6_0_cry_20_RNO_cZ.INIT=4'h6;
  LUT3 un9_6_0_cry_22_RNO_cZ(.I0(ZFF_Y1[5:5]),.I1(un9_11[22:22]),.I2(un9_11[26:26]),.O(un9_6_0_cry_22_RNO));
defparam un9_6_0_cry_22_RNO_cZ.INIT=8'h96;
  LUT3 un9_6_0_cry_23_RNO_cZ(.I0(un9_11[23:23]),.I1(ZFF_Y1[6:6]),.I2(ZFF_Y1[15:15]),.O(un9_6_0_cry_23_RNO));
defparam un9_6_0_cry_23_RNO_cZ.INIT=8'h96;
  LUT3 un9_6_0_cry_24_RNO_cZ(.I0(ZFF_Y1[7:7]),.I1(ZFF_Y1[16:16]),.I2(un9_11[24:24]),.O(un9_6_0_cry_24_RNO));
defparam un9_6_0_cry_24_RNO_cZ.INIT=8'h96;
  LUT3 un9_6_0_cry_25_RNO_cZ(.I0(ZFF_Y1[8:8]),.I1(un9_11[25:25]),.I2(ZFF_Y1[15:15]),.O(un9_6_0_cry_25_RNO));
defparam un9_6_0_cry_25_RNO_cZ.INIT=8'h96;
  LUT3 un9_6_0_cry_26_RNO_cZ(.I0(ZFF_Y1[9:9]),.I1(ZFF_Y1[16:16]),.I2(un9_11[26:26]),.O(un9_6_0_cry_26_RNO));
defparam un9_6_0_cry_26_RNO_cZ.INIT=8'h96;
  LUT3 un9_6_0_cry_28_RNO_cZ(.I0(un9_11[23:23]),.I1(ZFF_Y1[17:17]),.I2(un9_11[28:28]),.O(un9_6_0_cry_28_RNO));
defparam un9_6_0_cry_28_RNO_cZ.INIT=8'h96;
  LUT5 un9_11_s_8_RNIB86B1(.I0(ZFF_Y1_17_rep1),.I1(un9_11[23:23]),.I2(un9_11[24:24]),.I3(un9_11[29:29]),.I4(un9_11[28:28]),.O(un9_6_0_axb_29));
defparam un9_11_s_8_RNIB86B1.INIT=32'hE11E8778;
  LUT3 un9_6_0_cry_29_RNO_cZ(.I0(ZFF_Y1_17_rep1),.I1(un9_11[23:23]),.I2(un9_11[28:28]),.O(un9_6_0_cry_29_RNO));
defparam un9_6_0_cry_29_RNO_cZ.INIT=8'hE8;
  LUT5 un9_11_s_8_RNIHEPO1(.I0(un9_11[24:24]),.I1(un9_11[25:25]),.I2(ZFF_Y1[17:17]),.I3(un9_11[29:29]),.I4(un9_11[30:30]),.O(un9_6_0_axb_30));
defparam un9_11_s_8_RNIHEPO1.INIT=32'h69C3963C;
  LUT2 un9_6_0_cry_30_RNO_cZ(.I0(un9_11[24:24]),.I1(un9_11[29:29]),.O(un9_6_0_cry_30_RNO));
defparam un9_6_0_cry_30_RNO_cZ.INIT=4'h8;
  LUT5 un9_11_s_9_RNISG4V1(.I0(un9_11[25:25]),.I1(ZFF_Y1[17:17]),.I2(un9_11[26:26]),.I3(un9_11[30:30]),.I4(un9_11[31:31]),.O(un9_6_0_axb_31));
defparam un9_11_s_9_RNISG4V1.INIT=32'hE1871E78;
  LUT3 un9_6_0_cry_31_RNO_cZ(.I0(un9_11[25:25]),.I1(ZFF_Y1[17:17]),.I2(un9_11[30:30]),.O(un9_6_0_cry_31_RNO));
defparam un9_6_0_cry_31_RNO_cZ.INIT=8'hE8;
  LUT2 un9_6_0_cry_32_RNO_cZ(.I0(un9_11[26:26]),.I1(un9_11[31:31]),.O(un9_6_0_cry_32_RNO));
defparam un9_6_0_cry_32_RNO_cZ.INIT=4'h8;
  LUT2 un9_6_0_cry_33_RNO_cZ(.I0(ZFF_Y1[15:15]),.I1(un9_11[32:32]),.O(un9_6_0_cry_33_RNO));
defparam un9_6_0_cry_33_RNO_cZ.INIT=4'h8;
  LUT2 un9_6_0_cry_34_RNO_cZ(.I0(ZFF_Y1[16:16]),.I1(un9_11[33:33]),.O(un9_6_0_cry_34_RNO));
defparam un9_6_0_cry_34_RNO_cZ.INIT=4'h8;
  LUT2 un9_6_0_cry_35_RNO_cZ(.I0(ZFF_Y1[17:17]),.I1(un9_11[34:34]),.O(un9_6_0_cry_35_RNO));
defparam un9_6_0_cry_35_RNO_cZ.INIT=4'h8;
  LUT2 un9_6_0_cry_36_RNO_cZ(.I0(ZFF_Y1[17:17]),.I1(un9_11[35:35]),.O(un9_6_0_cry_36_RNO));
defparam un9_6_0_cry_36_RNO_cZ.INIT=4'h8;
  LUT2 un9_8_cry_6_RNO_cZ(.I0(un9_8_fast[6:6]),.I1(ZFF_Y1_fast[8:8]),.O(un9_8_cry_6_RNO));
defparam un9_8_cry_6_RNO_cZ.INIT=4'h8;
  LUT3 un9_8_cry_7_RNO_cZ(.I0(un9_8_fast[6:6]),.I1(ZFF_Y1_fast[5:5]),.I2(un9_11_fast[25:25]),.O(un9_8_cry_7_RNO));
defparam un9_8_cry_7_RNO_cZ.INIT=8'h96;
  LUT3 un9_8_cry_8_RNO_cZ(.I0(un9_8_7_rep1),.I1(un9_11_26_rep1),.I2(ZFF_Y1_6_rep1),.O(un9_8_cry_8_RNO));
defparam un9_8_cry_8_RNO_cZ.INIT=8'h96;
  LUT3 un9_8_cry_9_RNO_cZ(.I0(ZFF_Y1_9_rep1),.I1(ZFF_Y1_15_rep1),.I2(ZFF_Y1[3:3]),.O(un9_8_cry_9_RNO));
defparam un9_8_cry_9_RNO_cZ.INIT=8'h96;
  LUT3 un9_8_cry_10_RNO_cZ(.I0(un9_11_22_rep1),.I1(ZFF_Y1[4:4]),.I2(ZFF_Y1_16_rep1),.O(un9_8_cry_10_RNO));
defparam un9_8_cry_10_RNO_cZ.INIT=8'h96;
  LUT3 un9_8_cry_11_RNO_cZ(.I0(ZFF_Y1_9_rep1),.I1(un9_11_26_rep1),.I2(ZFF_Y1[5:5]),.O(un9_8_cry_11_RNO));
defparam un9_8_cry_11_RNO_cZ.INIT=8'h69;
  LUT3 un9_8_cry_12_RNO_cZ(.I0(ZFF_Y1_17_rep1),.I1(ZFF_Y1_6_rep1),.I2(un9_11_24_rep1),.O(un9_8_cry_12_RNO));
defparam un9_8_cry_12_RNO_cZ.INIT=8'h96;
  LUT3 un9_8_cry_13_RNO_cZ(.I0(ZFF_Y1_fast[17:17]),.I1(ZFF_Y1_fast[7:7]),.I2(un9_10_8_rep1),.O(un9_8_cry_13_RNO));
defparam un9_8_cry_13_RNO_cZ.INIT=8'h96;
  LUT3 un9_8_cry_17_RNO_cZ(.I0(ZFF_Y1_17_rep1),.I1(un9_11_fast[23:23]),.I2(ZFF_Y1_4_rep1),.O(un9_8_cry_17_RNO));
defparam un9_8_cry_17_RNO_cZ.INIT=8'h96;
  LUT2 un9_8_cry_21_RNO_cZ(.I0(ZFF_Y1[7:7]),.I1(un9_11[26:26]),.O(un9_8_cry_21_RNO));
defparam un9_8_cry_21_RNO_cZ.INIT=4'hB;
  LUT2 un9_8_cry_22_RNO_cZ(.I0(ZFF_Y1[8:8]),.I1(ZFF_Y1_15_rep1),.O(un9_8_cry_22_RNO));
defparam un9_8_cry_22_RNO_cZ.INIT=4'h2;
  LUT2 un9_8_cry_23_RNO_cZ(.I0(ZFF_Y1[9:9]),.I1(ZFF_Y1_16_rep1),.O(un9_8_cry_23_RNO));
defparam un9_8_cry_23_RNO_cZ.INIT=4'h2;
  LUT5 desc482(.I0(ZFF_Y1_fast[9:9]),.I1(un9_8_7_rep1),.I2(ZFF_Y1_3_rep1),.I3(ZFF_Y1_7_rep1),.I4(ZFF_Y1_4_rep1),.O(un9_10_axb_3));
defparam desc482.INIT=32'hE11E8778;
  LUT3 un9_10_cry_3_RNO_cZ(.I0(ZFF_Y1_fast[9:9]),.I1(un9_8_7_rep1),.I2(ZFF_Y1_4_rep1),.O(un9_10_cry_3_RNO));
defparam un9_10_cry_3_RNO_cZ.INIT=8'hE8;
  LUT2 un9_10_cry_4_RNO_cZ(.I0(ZFF_Y1_3_rep1),.I1(ZFF_Y1_7_rep1),.O(un9_10_cry_4_RNO));
defparam un9_10_cry_4_RNO_cZ.INIT=4'h8;
  LUT5 desc483(.I0(un9_11_fast[24:24]),.I1(ZFF_Y1_fast[8:8]),.I2(ZFF_Y1_5_rep1),.I3(ZFF_Y1_7_rep1),.I4(ZFF_Y1_4_rep1),.O(un9_10_axb_5));
defparam desc483.INIT=32'h6996A55A;
  LUT2 un9_10_cry_5_RNO_cZ(.I0(ZFF_Y1_fast[8:8]),.I1(ZFF_Y1_4_rep1),.O(un9_10_cry_5_RNO));
defparam un9_10_cry_5_RNO_cZ.INIT=4'h8;
  LUT3 un9_10_cry_6_RNO_cZ(.I0(ZFF_Y1[6:6]),.I1(ZFF_Y1[8:8]),.I2(un9_11[25:25]),.O(un9_10_cry_6_RNO));
defparam un9_10_cry_6_RNO_cZ.INIT=8'h96;
  LUT5 desc484(.I0(un9_11_fast[25:25]),.I1(ZFF_Y1_6_rep1),.I2(ZFF_Y1_fast[8:8]),.I3(ZFF_Y1_7_rep1),.I4(un9_10_8_rep1),.O(un9_10_axb_7));
defparam desc484.INIT=32'hE81717E8;
  LUT3 un9_10_cry_7_RNO_cZ(.I0(un9_11_fast[25:25]),.I1(ZFF_Y1_6_rep1),.I2(ZFF_Y1_fast[8:8]),.O(un9_10_cry_7_RNO));
defparam un9_10_cry_7_RNO_cZ.INIT=8'hE8;
  LUT5 ZFF_Y1_10_rep1_RNIP55H1(.I0(un9_11_22_rep1),.I1(un9_8_6_rep1),.I2(ZFF_Y1_fast[8:8]),.I3(ZFF_Y1_7_rep1),.I4(un9_10_8_rep1),.O(un9_10_axb_8));
defparam ZFF_Y1_10_rep1_RNIP55H1.INIT=32'h69969696;
  LUT2 un9_10_cry_8_RNO_cZ(.I0(ZFF_Y1_7_rep1),.I1(un9_10_8_rep1),.O(un9_10_cry_8_RNO));
defparam un9_10_cry_8_RNO_cZ.INIT=4'h8;
  LUT3 un9_10_cry_9_RNO_cZ(.I0(un9_11[23:23]),.I1(un9_11[25:25]),.I2(un9_8[7:7]),.O(un9_10_cry_9_RNO));
defparam un9_10_cry_9_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_10_RNO_cZ(.I0(un9_11[24:24]),.I1(ZFF_Y1[3:3]),.I2(un9_10[8:8]),.O(un9_10_cry_10_RNO));
defparam un9_10_cry_10_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_11_RNO_cZ(.I0(un9_8[6:6]),.I1(ZFF_Y1[4:4]),.I2(un9_11[25:25]),.O(un9_10_cry_11_RNO));
defparam un9_10_cry_11_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_12_RNO_cZ(.I0(ZFF_Y1[5:5]),.I1(un9_8[7:7]),.I2(un9_11[26:26]),.O(un9_10_cry_12_RNO));
defparam un9_10_cry_12_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_13_RNO_cZ(.I0(ZFF_Y1[6:6]),.I1(ZFF_Y1[3:3]),.I2(un9_10[8:8]),.O(un9_10_cry_13_RNO));
defparam un9_10_cry_13_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_14_RNO_cZ(.I0(un9_8[6:6]),.I1(ZFF_Y1[7:7]),.I2(ZFF_Y1[4:4]),.O(un9_10_cry_14_RNO));
defparam un9_10_cry_14_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_15_RNO_cZ(.I0(ZFF_Y1[5:5]),.I1(ZFF_Y1[8:8]),.I2(un9_8[7:7]),.O(un9_10_cry_15_RNO));
defparam un9_10_cry_15_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_16_RNO_cZ(.I0(ZFF_Y1[9:9]),.I1(ZFF_Y1[6:6]),.I2(ZFF_Y1[3:3]),.O(un9_10_cry_16_RNO));
defparam un9_10_cry_16_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_17_RNO_cZ(.I0(ZFF_Y1[7:7]),.I1(ZFF_Y1[4:4]),.I2(un9_11[22:22]),.O(un9_10_cry_17_RNO));
defparam un9_10_cry_17_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_18_RNO_cZ(.I0(un9_11[23:23]),.I1(ZFF_Y1[5:5]),.I2(ZFF_Y1[8:8]),.O(un9_10_cry_18_RNO));
defparam un9_10_cry_18_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_19_RNO_cZ(.I0(ZFF_Y1[9:9]),.I1(ZFF_Y1[6:6]),.I2(un9_11[24:24]),.O(un9_10_cry_19_RNO));
defparam un9_10_cry_19_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_20_RNO_cZ(.I0(ZFF_Y1[7:7]),.I1(un9_11[25:25]),.I2(un9_11[22:22]),.O(un9_10_cry_20_RNO));
defparam un9_10_cry_20_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_21_RNO_cZ(.I0(un9_11[23:23]),.I1(ZFF_Y1[8:8]),.I2(un9_11[26:26]),.O(un9_10_cry_21_RNO));
defparam un9_10_cry_21_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_22_RNO_cZ(.I0(ZFF_Y1[9:9]),.I1(un9_11[24:24]),.I2(ZFF_Y1[15:15]),.O(un9_10_cry_22_RNO));
defparam un9_10_cry_22_RNO_cZ.INIT=8'h96;
  LUT3 un9_10_cry_23_RNO_cZ(.I0(ZFF_Y1[16:16]),.I1(un9_11[25:25]),.I2(un9_11[22:22]),.O(un9_10_cry_23_RNO));
defparam un9_10_cry_23_RNO_cZ.INIT=8'h96;
  LUT5 ZFF_Y1_11_rep1_RNIGK1E1(.I0(un9_11_23_rep1),.I1(un9_11_25_rep1),.I2(ZFF_Y1_16_rep1),.I3(un9_11[22:22]),.I4(un9_11[26:26]),.O(un9_10_axb_24));
defparam ZFF_Y1_11_rep1_RNIGK1E1.INIT=32'hA995566A;
  LUT3 un9_10_cry_24_RNO_cZ(.I0(un9_11_25_rep1),.I1(ZFF_Y1_16_rep1),.I2(un9_11[22:22]),.O(un9_10_cry_24_RNO));
defparam un9_10_cry_24_RNO_cZ.INIT=8'hE8;
  LUT2 un9_10_cry_25_RNO_cZ(.I0(un9_11[23:23]),.I1(un9_11[26:26]),.O(un9_10_cry_25_RNO));
defparam un9_10_cry_25_RNO_cZ.INIT=4'h8;
  LUT2 un9_10_cry_26_RNO_cZ(.I0(un9_11[24:24]),.I1(ZFF_Y1[15:15]),.O(un9_10_cry_26_RNO));
defparam un9_10_cry_26_RNO_cZ.INIT=4'h8;
  LUT2 un9_10_cry_27_RNO_cZ(.I0(ZFF_Y1[16:16]),.I1(un9_11[25:25]),.O(un9_10_cry_27_RNO));
defparam un9_10_cry_27_RNO_cZ.INIT=4'h8;
  LUT2 un10_cry_29_RNO_cZ(.I0(un10_8[35:35]),.I1(un10_6[35:35]),.O(un10_cry_29_RNO));
defparam un10_cry_29_RNO_cZ.INIT=4'h6;
  LUT2 un10_cry_30_RNO_cZ(.I0(un10_8[35:35]),.I1(un10_6[35:35]),.O(un10_cry_30_RNO));
defparam un10_cry_30_RNO_cZ.INIT=4'h8;
  LUT2 un10_cry_31_RNO_cZ(.I0(un10_8[36:36]),.I1(un10_6[36:36]),.O(un10_cry_31_RNO));
defparam un10_cry_31_RNO_cZ.INIT=4'hE;
  LUT5 desc485(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[0:0]),.I2(ZFF_Y2[2:2]),.I3(ZFF_Y2[1:1]),.I4(ZFF_Y2[9:9]),.O(un10_6[9:9]));
defparam desc485.INIT=32'hD42B2BD4;
  LUT3 un10_6_cry_0_RNO_cZ(.I0(ZFF_Y2_fast[8:8]),.I1(ZFF_Y2[0:0]),.I2(ZFF_Y2[2:2]),.O(un10_6_cry_0_RNO));
defparam un10_6_cry_0_RNO_cZ.INIT=8'h2B;
  LUT2 un10_6_cry_1_RNO_cZ(.I0(ZFF_Y2[1:1]),.I1(ZFF_Y2[9:9]),.O(un10_6_cry_1_RNO));
defparam un10_6_cry_1_RNO_cZ.INIT=4'h4;
  LUT2 un10_6_cry_2_RNO_cZ(.I0(ZFF_Y2[2:2]),.I1(ZFF_Y2[10:10]),.O(un10_6_cry_2_RNO));
defparam un10_6_cry_2_RNO_cZ.INIT=4'h4;
  LUT5 desc486(.I0(ZFF_Y2[4:4]),.I1(ZFF_Y2[0:0]),.I2(ZFF_Y2[3:3]),.I3(ZFF_Y2[12:12]),.I4(ZFF_Y2[11:11]),.O(un10_6_axb_3));
defparam desc486.INIT=32'h69966699;
  LUT2 un10_6_cry_3_RNO_cZ(.I0(ZFF_Y2[3:3]),.I1(ZFF_Y2[11:11]),.O(un10_6_cry_3_RNO));
defparam un10_6_cry_3_RNO_cZ.INIT=4'h4;
  LUT3 un10_6_cry_4_RNO_cZ(.I0(ZFF_Y2[5:5]),.I1(ZFF_Y2[1:1]),.I2(ZFF_Y2[13:13]),.O(un10_6_cry_4_RNO));
defparam un10_6_cry_4_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_5_RNO_cZ(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[0:0]),.I2(ZFF_Y2[2:2]),.O(un10_6_cry_5_RNO));
defparam un10_6_cry_5_RNO_cZ.INIT=8'h96;
  LUT3 un10_6_cry_6_RNO_cZ(.I0(ZFF_Y2[3:3]),.I1(ZFF_Y2[1:1]),.I2(ZFF_Y2[15:15]),.O(un10_6_cry_6_RNO));
defparam un10_6_cry_6_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_7_RNO_cZ(.I0(ZFF_Y2[4:4]),.I1(ZFF_Y2[2:2]),.I2(ZFF_Y2[16:16]),.O(un10_6_cry_7_RNO));
defparam un10_6_cry_7_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_8_RNO_cZ(.I0(ZFF_Y2[5:5]),.I1(ZFF_Y2[3:3]),.I2(ZFF_Y2[9:9]),.O(un10_6_cry_8_RNO));
defparam un10_6_cry_8_RNO_cZ.INIT=8'h96;
  LUT3 un10_6_cry_9_RNO_cZ(.I0(ZFF_Y2_6_rep1),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[0:0]),.O(un10_6_cry_9_RNO));
defparam un10_6_cry_9_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_10_RNO_cZ(.I0(ZFF_Y2_7_rep1),.I1(ZFF_Y2[5:5]),.I2(ZFF_Y2[1:1]),.O(un10_6_cry_10_RNO));
defparam un10_6_cry_10_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_11_RNO_cZ(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[6:6]),.I2(ZFF_Y2[2:2]),.O(un10_6_cry_11_RNO));
defparam un10_6_cry_11_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_12_RNO_cZ(.I0(ZFF_Y2_7_rep1),.I1(ZFF_Y2[3:3]),.I2(ZFF_Y2[9:9]),.O(un10_6_cry_12_RNO));
defparam un10_6_cry_12_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_13_RNO_cZ(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[4:4]),.I2(ZFF_Y2[10:10]),.O(un10_6_cry_13_RNO));
defparam un10_6_cry_13_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_14_RNO_cZ(.I0(ZFF_Y2[5:5]),.I1(ZFF_Y2[11:11]),.I2(ZFF_Y2[9:9]),.O(un10_6_cry_14_RNO));
defparam un10_6_cry_14_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_15_RNO_cZ(.I0(ZFF_Y2[6:6]),.I1(ZFF_Y2[12:12]),.I2(ZFF_Y2[10:10]),.O(un10_6_cry_15_RNO));
defparam un10_6_cry_15_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_16_RNO_cZ(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[11:11]),.I2(ZFF_Y2[13:13]),.O(un10_6_cry_16_RNO));
defparam un10_6_cry_16_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_17_RNO_cZ(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[14:14]),.I2(ZFF_Y2[12:12]),.O(un10_6_cry_17_RNO));
defparam un10_6_cry_17_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_18_RNO_cZ(.I0(ZFF_Y2[13:13]),.I1(ZFF_Y2[15:15]),.I2(ZFF_Y2[9:9]),.O(un10_6_cry_18_RNO));
defparam un10_6_cry_18_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_19_RNO_cZ(.I0(ZFF_Y2[14:14]),.I1(ZFF_Y2[10:10]),.I2(ZFF_Y2[16:16]),.O(un10_6_cry_19_RNO));
defparam un10_6_cry_19_RNO_cZ.INIT=8'h69;
  LUT3 un10_6_cry_20_RNO_cZ(.I0(ZFF_Y2_14_rep1),.I1(ZFF_Y2[10:10]),.I2(ZFF_Y2[16:16]),.O(un10_6_cry_20_RNO));
defparam un10_6_cry_20_RNO_cZ.INIT=8'hD4;
  LUT2 un10_6_cry_21_RNO_cZ(.I0(ZFF_Y2[11:11]),.I1(ZFF_Y2[15:15]),.O(un10_6_cry_21_RNO));
defparam un10_6_cry_21_RNO_cZ.INIT=4'h2;
  LUT2 un10_6_cry_22_RNO_cZ(.I0(ZFF_Y2[12:12]),.I1(ZFF_Y2[16:16]),.O(un10_6_cry_22_RNO));
defparam un10_6_cry_22_RNO_cZ.INIT=4'h2;
  LUT2 un10_6_cry_23_RNO_cZ(.I0(ZFF_Y2[13:13]),.I1(ZFF_Y2[17:17]),.O(un10_6_cry_23_RNO));
defparam un10_6_cry_23_RNO_cZ.INIT=4'h2;
  LUT2 un10_6_cry_24_RNO(.I0(ZFF_Y2[14:14]),.I1(ZFF_Y2[17:17]),.O(un10_8_34));
defparam un10_6_cry_24_RNO.INIT=4'h2;
  LUT2 un10_6_cry_25_RNO(.I0(ZFF_Y2[15:15]),.I1(ZFF_Y2[17:17]),.O(un10_8_37));
defparam un10_6_cry_25_RNO.INIT=4'h2;
  LUT2 un10_6_cry_26_RNO(.I0(ZFF_Y2[16:16]),.I1(ZFF_Y2[17:17]),.O(un10_8_40));
defparam un10_6_cry_26_RNO.INIT=4'h2;
  LUT5 un8_0_8_s_18_RNITBHC1(.I0(un8_0_6[28:28]),.I1(un8_0_8[28:28]),.I2(un8_0_9[28:28]),.I3(un8_0_8[29:29]),.I4(un8_0_9[29:29]),.O(un8_0_0_axb_29));
defparam un8_0_8_s_18_RNITBHC1.INIT=32'hE81717E8;
  LUT2 un8_0_0_cry_29_RNO_cZ(.I0(un8_0_8[29:29]),.I1(un8_0_9[29:29]),.O(un8_0_0_cry_29_RNO));
defparam un8_0_0_cry_29_RNO_cZ.INIT=4'h6;
  LUT2 un8_0_0_cry_30_RNO_cZ(.I0(un8_0_8[29:29]),.I1(un8_0_9[29:29]),.O(un8_0_0_cry_30_RNO));
defparam un8_0_0_cry_30_RNO_cZ.INIT=4'h8;
  LUT2 un8_0_0_cry_31_RNO_cZ(.I0(un8_0_8[30:30]),.I1(un8_0_9[30:30]),.O(un8_0_0_cry_31_RNO));
defparam un8_0_0_cry_31_RNO_cZ.INIT=4'h8;
  LUT2 un8_0_0_cry_32_RNO_cZ(.I0(un8_0_8[31:31]),.I1(un8_0_9[31:31]),.O(un8_0_0_cry_32_RNO));
defparam un8_0_0_cry_32_RNO_cZ.INIT=4'h8;
  LUT2 un8_0_0_cry_33_RNO_cZ(.I0(un8_0_8[32:32]),.I1(un8_0_9[32:32]),.O(un8_0_0_cry_33_RNO));
defparam un8_0_0_cry_33_RNO_cZ.INIT=4'h8;
  LUT2 un8_0_0_cry_34_RNO_cZ(.I0(un8_0_8[33:33]),.I1(un8_0_9[33:33]),.O(un8_0_0_cry_34_RNO));
defparam un8_0_0_cry_34_RNO_cZ.INIT=4'h8;
  LUT2 un8_0_0_cry_35_RNO_cZ(.I0(un8_0_8[34:34]),.I1(un8_0_9[34:34]),.O(un8_0_0_cry_35_RNO));
defparam un8_0_0_cry_35_RNO_cZ.INIT=4'h8;
  LUT2 un8_0_0_cry_36_RNO_cZ(.I0(un8_0_8[35:35]),.I1(un8_0_9[35:35]),.O(un8_0_0_cry_36_RNO));
defparam un8_0_0_cry_36_RNO_cZ.INIT=4'h8;
  LUT5 ZFF_X2_2_rep1_RNI2DGC1(.I0(ZFF_X2_2_rep1),.I1(ZFF_X2_3_rep1),.I2(ZFF_X2[4:4]),.I3(ZFF_X2[9:9]),.I4(ZFF_X2[1:1]),.O(un8_0_6_axb_4));
defparam ZFF_X2_2_rep1_RNI2DGC1.INIT=32'h96695AA5;
  LUT2 un8_0_6_cry_4_RNO_cZ(.I0(ZFF_X2_3_rep1),.I1(ZFF_X2[1:1]),.O(un8_0_6_cry_4_RNO));
defparam un8_0_6_cry_4_RNO_cZ.INIT=4'h8;
  LUT3 un8_0_6_cry_5_RNO_cZ(.I0(ZFF_X2[0:0]),.I1(ZFF_X2[10:10]),.I2(ZFF_X2[5:5]),.O(un8_0_6_cry_5_RNO));
defparam un8_0_6_cry_5_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_6_RNO_cZ(.I0(ZFF_X2[6:6]),.I1(ZFF_X2[1:1]),.I2(ZFF_X2[11:11]),.O(un8_0_6_cry_6_RNO));
defparam un8_0_6_cry_6_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_7_RNO_cZ(.I0(ZFF_X2[2:2]),.I1(ZFF_X2[0:0]),.I2(ZFF_X2[12:12]),.O(un8_0_6_cry_7_RNO));
defparam un8_0_6_cry_7_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_8_RNO_cZ(.I0(ZFF_X2[3:3]),.I1(ZFF_X2[1:1]),.I2(ZFF_X2[13:13]),.O(un8_0_6_cry_8_RNO));
defparam un8_0_6_cry_8_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_9_RNO_cZ(.I0(ZFF_X2[14:14]),.I1(ZFF_X2[2:2]),.I2(ZFF_X2[4:4]),.O(un8_0_6_cry_9_RNO));
defparam un8_0_6_cry_9_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_10_RNO_cZ(.I0(ZFF_X2[3:3]),.I1(ZFF_X2[5:5]),.I2(ZFF_X2[15:15]),.O(un8_0_6_cry_10_RNO));
defparam un8_0_6_cry_10_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_11_RNO_cZ(.I0(ZFF_X2[4:4]),.I1(ZFF_X2[6:6]),.I2(ZFF_X2[16:16]),.O(un8_0_6_cry_11_RNO));
defparam un8_0_6_cry_11_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_12_RNO_cZ(.I0(ZFF_X2[5:5]),.I1(ZFF_X2[7:7]),.I2(ZFF_X2_fast[16:16]),.O(un8_0_6_cry_12_RNO));
defparam un8_0_6_cry_12_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_13_RNO_cZ(.I0(ZFF_X2[6:6]),.I1(ZFF_X2[8:8]),.I2(ZFF_X2_fast[16:16]),.O(un8_0_6_cry_13_RNO));
defparam un8_0_6_cry_13_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_14_RNO_cZ(.I0(ZFF_X2[9:9]),.I1(ZFF_X2[7:7]),.I2(ZFF_X2_fast[16:16]),.O(un8_0_6_cry_14_RNO));
defparam un8_0_6_cry_14_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_15_RNO_cZ(.I0(ZFF_X2[10:10]),.I1(ZFF_X2[8:8]),.I2(ZFF_X2_fast[16:16]),.O(un8_0_6_cry_15_RNO));
defparam un8_0_6_cry_15_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_6_cry_16_RNO_cZ(.I0(ZFF_X2[10:10]),.I1(ZFF_X2[16:16]),.I2(ZFF_X2[8:8]),.O(un8_0_6_cry_16_RNO));
defparam un8_0_6_cry_16_RNO_cZ.INIT=8'hB2;
  LUT3 un8_0_6_cry_17_RNO_cZ(.I0(ZFF_X2[10:10]),.I1(ZFF_X2[15:15]),.I2(ZFF_X2[12:12]),.O(un8_0_6_cry_17_RNO));
defparam un8_0_6_cry_17_RNO_cZ.INIT=8'h96;
  LUT3 un8_0_6_cry_18_RNO_cZ(.I0(ZFF_X2[15:15]),.I1(ZFF_X2[13:13]),.I2(ZFF_X2[11:11]),.O(un8_0_6_cry_18_RNO));
defparam un8_0_6_cry_18_RNO_cZ.INIT=8'h96;
  LUT5 ZFF_X2_14_rep1_RNILO071(.I0(ZFF_X2_14_rep1),.I1(ZFF_X2[15:15]),.I2(ZFF_X2[12:12]),.I3(ZFF_X2[13:13]),.I4(ZFF_X2[11:11]),.O(un8_0_6_axb_19));
defparam ZFF_X2_14_rep1_RNILO071.INIT=32'hA596965A;
  LUT3 un8_0_6_cry_19_RNO_cZ(.I0(ZFF_X2[15:15]),.I1(ZFF_X2[13:13]),.I2(ZFF_X2[11:11]),.O(un8_0_6_cry_19_RNO));
defparam un8_0_6_cry_19_RNO_cZ.INIT=8'hE8;
  LUT2 un8_0_6_cry_20_RNO_cZ(.I0(ZFF_X2_14_rep1),.I1(ZFF_X2[12:12]),.O(un8_0_6_cry_20_RNO));
defparam un8_0_6_cry_20_RNO_cZ.INIT=4'h8;
  LUT2 un8_0_6_cry_21_RNO(.I0(ZFF_X2[15:15]),.I1(ZFF_X2[13:13]),.O(un8_0_6_43));
defparam un8_0_6_cry_21_RNO.INIT=4'h8;
  LUT2 desc487(.I0(ZFF_X1_fast[0:0]),.I1(ZFF_X1_fast[3:3]),.O(un7_0_8[9:9]));
defparam desc487.INIT=4'h6;
  LUT5 un7_0_10_s_15_RNIDDTA1(.I0(un7_0_6[33:33]),.I1(un7_0_10[33:33]),.I2(un7_0_8[33:33]),.I3(un7_0_10[34:34]),.I4(un7_0_8[34:34]),.O(un7_0_0_axb_34));
defparam un7_0_10_s_15_RNIDDTA1.INIT=32'hE81717E8;
  LUT2 un7_0_0_cry_34_RNO_cZ(.I0(un7_0_10[34:34]),.I1(un7_0_8[34:34]),.O(un7_0_0_cry_34_RNO));
defparam un7_0_0_cry_34_RNO_cZ.INIT=4'h6;
  LUT2 un7_0_0_cry_35_RNO_cZ(.I0(un7_0_10[34:34]),.I1(un7_0_8[34:34]),.O(un7_0_0_cry_35_RNO));
defparam un7_0_0_cry_35_RNO_cZ.INIT=4'h8;
  LUT2 un7_0_0_cry_36_RNO_cZ(.I0(un7_0_10[35:35]),.I1(un7_0_8[35:35]),.O(un7_0_0_cry_36_RNO));
defparam un7_0_0_cry_36_RNO_cZ.INIT=4'h8;
  LUT2 un7_0_0_cry_37_RNO_cZ(.I0(un7_0_10[36:36]),.I1(un7_0_8[36:36]),.O(un7_0_0_cry_37_RNO));
defparam un7_0_0_cry_37_RNO_cZ.INIT=4'h8;
  LUT5 un7_0_10_s_20_RNI6UHP(.I0(ZFF_X1[16:16]),.I1(un7_0_8[38:38]),.I2(un7_0_10[38:38]),.I3(un7_0_10[37:37]),.I4(un7_0_8[37:37]),.O(un7_0_0_axb_38));
defparam un7_0_10_s_20_RNI6UHP.INIT=32'h69969696;
  LUT2 un7_0_0_cry_38_RNO_cZ(.I0(un7_0_10[37:37]),.I1(un7_0_8[37:37]),.O(un7_0_0_cry_38_RNO));
defparam un7_0_0_cry_38_RNO_cZ.INIT=4'h8;
  LUT2 un7_0_0_cry_39_RNO_cZ(.I0(ZFF_X1[16:16]),.I1(un7_0_10[39:39]),.O(un7_0_0_cry_39_RNO));
defparam un7_0_0_cry_39_RNO_cZ.INIT=4'h6;
  LUT2 un7_0_0_cry_40_RNO_cZ(.I0(ZFF_X1[16:16]),.I1(un7_0_10[39:39]),.O(un7_0_0_cry_40_RNO));
defparam un7_0_0_cry_40_RNO_cZ.INIT=4'h8;
  LUT2 un7_0_0_cry_41_RNO_cZ(.I0(ZFF_X1[16:16]),.I1(un7_0_10[40:40]),.O(un7_0_0_cry_41_RNO));
defparam un7_0_0_cry_41_RNO_cZ.INIT=4'h8;
  LUT5 desc488(.I0(ZFF_X1_fast[0:0]),.I1(ZFF_X1_fast[7:7]),.I2(ZFF_X1_fast[1:1]),.I3(ZFF_X1_fast[3:3]),.I4(ZFF_X1_fast[4:4]),.O(un7_0_6_axb_4));
defparam desc488.INIT=32'h963C69C3;
  LUT2 un7_0_6_cry_4_RNO_cZ(.I0(ZFF_X1_fast[0:0]),.I1(ZFF_X1_fast[3:3]),.O(un7_0_6_cry_4_RNO));
defparam un7_0_6_cry_4_RNO_cZ.INIT=4'h8;
  LUT5 desc489(.I0(ZFF_X1_fast[7:7]),.I1(ZFF_X1_fast[1:1]),.I2(ZFF_X1_fast[8:8]),.I3(ZFF_X1_fast[2:2]),.I4(ZFF_X1_fast[4:4]),.O(un7_0_6_axb_5));
defparam desc489.INIT=32'h2DD2B44B;
  LUT3 un7_0_6_cry_5_RNO_cZ(.I0(ZFF_X1_fast[7:7]),.I1(ZFF_X1_fast[1:1]),.I2(ZFF_X1_fast[4:4]),.O(un7_0_6_cry_5_RNO));
defparam un7_0_6_cry_5_RNO_cZ.INIT=8'hD4;
  LUT2 un7_0_6_cry_6_RNO_cZ(.I0(ZFF_X1_fast[8:8]),.I1(ZFF_X1_fast[2:2]),.O(un7_0_6_cry_6_RNO));
defparam un7_0_6_cry_6_RNO_cZ.INIT=4'h4;
  LUT2 un7_0_6_cry_7_RNO(.I0(ZFF_X1_fast[6:6]),.I1(ZFF_X1_9_rep1),.O(un7_0_10_14));
defparam un7_0_6_cry_7_RNO.INIT=4'h2;
  LUT2 un7_0_6_cry_8_RNO_cZ(.I0(ZFF_X1_fast[10:10]),.I1(ZFF_X1_0_rep1),.O(un7_0_6_cry_8_RNO));
defparam un7_0_6_cry_8_RNO_cZ.INIT=4'h4;
  LUT2 un7_0_6_cry_9_RNO_cZ(.I0(ZFF_X1_fast[11:11]),.I1(ZFF_X1_1_rep1),.O(un7_0_6_cry_9_RNO));
defparam un7_0_6_cry_9_RNO_cZ.INIT=4'h4;
  LUT3 un7_0_6_cry_10_RNO_cZ(.I0(ZFF_X1_fast[13:13]),.I1(ZFF_X1_fast[3:3]),.I2(ZFF_X1_fast[4:4]),.O(un7_0_6_cry_10_RNO));
defparam un7_0_6_cry_10_RNO_cZ.INIT=8'h69;
  LUT3 un7_0_6_cry_11_RNO_cZ(.I0(ZFF_X1_fast[8:8]),.I1(ZFF_X1_fast[4:4]),.I2(ZFF_X1_fast[14:14]),.O(un7_0_6_cry_11_RNO));
defparam un7_0_6_cry_11_RNO_cZ.INIT=8'h69;
  LUT3 un7_0_6_cry_12_RNO_cZ(.I0(ZFF_X1_5_rep1),.I1(ZFF_X1_9_rep1),.I2(ZFF_X1_15_rep1),.O(un7_0_6_cry_12_RNO));
defparam un7_0_6_cry_12_RNO_cZ.INIT=8'h69;
  LUT3 un7_0_6_cry_13_RNO_cZ(.I0(ZFF_X1_6_rep1),.I1(ZFF_X1_10_rep1),.I2(ZFF_X1_fast[16:16]),.O(un7_0_6_cry_13_RNO));
defparam un7_0_6_cry_13_RNO_cZ.INIT=8'h69;
  LUT3 un7_0_6_cry_14_RNO_cZ(.I0(ZFF_X1_0_rep1),.I1(ZFF_X1_7_rep1),.I2(ZFF_X1_fast[16:16]),.O(un7_0_6_cry_14_RNO));
defparam un7_0_6_cry_14_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_6_cry_15_RNO_cZ(.I0(ZFF_X1_1_rep1),.I1(ZFF_X1_8_rep1),.I2(ZFF_X1_fast[16:16]),.O(un7_0_6_cry_15_RNO));
defparam un7_0_6_cry_15_RNO_cZ.INIT=8'h96;
  LUT2 un7_0_6_cry_22_RNO_cZ(.I0(ZFF_X1_7_rep1),.I1(ZFF_X1[14:14]),.O(un7_0_6_cry_22_RNO));
defparam un7_0_6_cry_22_RNO_cZ.INIT=4'hD;
  LUT2 un7_0_6_cry_23_RNO_cZ(.I0(ZFF_X1_15_rep1),.I1(ZFF_X1_8_rep1),.O(un7_0_6_cry_23_RNO));
defparam un7_0_6_cry_23_RNO_cZ.INIT=4'h2;
  LUT3 un7_0_8_cry_6_RNO_cZ(.I0(ZFF_X1_6_rep1),.I1(ZFF_X1[3:3]),.I2(ZFF_X1[1:1]),.O(un7_0_8_cry_6_RNO));
defparam un7_0_8_cry_6_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_7_RNO_cZ(.I0(ZFF_X1_2_rep1),.I1(ZFF_X1_7_rep1),.I2(ZFF_X1[4:4]),.O(un7_0_8_cry_7_RNO));
defparam un7_0_8_cry_7_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_8_RNO_cZ(.I0(ZFF_X1[3:3]),.I1(ZFF_X1[5:5]),.I2(ZFF_X1[14:14]),.O(un7_0_8_cry_8_RNO));
defparam un7_0_8_cry_8_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_9_RNO_cZ(.I0(ZFF_X1_12_rep1),.I1(ZFF_X1[4:4]),.I2(ZFF_X1[6:6]),.O(un7_0_8_cry_9_RNO));
defparam un7_0_8_cry_9_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_10_RNO_cZ(.I0(ZFF_X1_13_rep1),.I1(ZFF_X1[5:5]),.I2(ZFF_X1[7:7]),.O(un7_0_8_cry_10_RNO));
defparam un7_0_8_cry_10_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_11_RNO_cZ(.I0(ZFF_X1_8_rep1),.I1(ZFF_X1[6:6]),.I2(ZFF_X1[14:14]),.O(un7_0_8_cry_11_RNO));
defparam un7_0_8_cry_11_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_12_RNO_cZ(.I0(ZFF_X1[15:15]),.I1(ZFF_X1[9:9]),.I2(ZFF_X1[7:7]),.O(un7_0_8_cry_12_RNO));
defparam un7_0_8_cry_12_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_13_RNO_cZ(.I0(ZFF_X1[0:0]),.I1(ZFF_X1[8:8]),.I2(ZFF_X1[10:10]),.O(un7_0_8_cry_13_RNO));
defparam un7_0_8_cry_13_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_14_RNO_cZ(.I0(ZFF_X1_11_rep1),.I1(ZFF_X1[1:1]),.I2(ZFF_X1[9:9]),.O(un7_0_8_cry_14_RNO));
defparam un7_0_8_cry_14_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_15_RNO_cZ(.I0(ZFF_X1_12_rep1),.I1(ZFF_X1[2:2]),.I2(ZFF_X1[10:10]),.O(un7_0_8_cry_15_RNO));
defparam un7_0_8_cry_15_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_16_RNO_cZ(.I0(ZFF_X1_11_rep1),.I1(ZFF_X1[3:3]),.I2(ZFF_X1[13:13]),.O(un7_0_8_cry_16_RNO));
defparam un7_0_8_cry_16_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_17_RNO_cZ(.I0(ZFF_X1[4:4]),.I1(ZFF_X1[12:12]),.I2(ZFF_X1[14:14]),.O(un7_0_8_cry_17_RNO));
defparam un7_0_8_cry_17_RNO_cZ.INIT=8'h96;
  LUT3 un7_0_8_cry_18_RNO_cZ(.I0(ZFF_X1[5:5]),.I1(ZFF_X1[13:13]),.I2(ZFF_X1[15:15]),.O(un7_0_8_cry_18_RNO));
defparam un7_0_8_cry_18_RNO_cZ.INIT=8'h96;
  LUT5 ZFF_X1_5_rep1_RNITSMV(.I0(ZFF_X1_5_rep1),.I1(ZFF_X1_6_rep1),.I2(ZFF_X1_13_rep1),.I3(ZFF_X1_15_rep1),.I4(ZFF_X1_fast[14:14]),.O(un7_0_8_axb_19));
defparam ZFF_X1_5_rep1_RNITSMV.INIT=32'hC993366C;
  LUT3 un7_0_8_cry_19_RNO_cZ(.I0(ZFF_X1_5_rep1),.I1(ZFF_X1_13_rep1),.I2(ZFF_X1_15_rep1),.O(un7_0_8_cry_19_RNO));
defparam un7_0_8_cry_19_RNO_cZ.INIT=8'hE8;
  LUT2 un7_0_8_cry_20_RNO(.I0(ZFF_X1_6_rep1),.I1(ZFF_X1_fast[14:14]),.O(un7_0_8_19));
defparam un7_0_8_cry_20_RNO.INIT=4'h8;
  LUT2 un7_0_8_cry_21_RNO(.I0(ZFF_X1[15:15]),.I1(ZFF_X1[7:7]),.O(un7_0_8_22));
defparam un7_0_8_cry_21_RNO.INIT=4'h8;
  LUT3 un6_0_8_cry_3_RNO_cZ(.I0(ZFF_X0_fast[6:6]),.I1(ZFF_X0_fast[8:8]),.I2(ZFF_X0_fast[5:5]),.O(un6_0_8_cry_3_RNO));
defparam un6_0_8_cry_3_RNO_cZ.INIT=8'h96;
  LUT3 un6_0_8_cry_4_RNO_cZ(.I0(ZFF_X0_fast[7:7]),.I1(ZFF_X0_fast[6:6]),.I2(ZFF_X0_fast[9:9]),.O(un6_0_8_cry_4_RNO));
defparam un6_0_8_cry_4_RNO_cZ.INIT=8'h96;
  LUT3 un6_0_8_cry_6_RNO_cZ(.I0(ZFF_X0_fast[1:1]),.I1(ZFF_X0_fast[11:11]),.I2(ZFF_X0_fast[9:9]),.O(un6_0_8_cry_6_RNO));
defparam un6_0_8_cry_6_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_8_cry_7_RNO_cZ(.I0(ZFF_X0_2_rep1),.I1(ZFF_X0_10_rep1),.I2(ZFF_X0_12_rep1),.O(un6_0_8_cry_7_RNO));
defparam un6_0_8_cry_7_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_8_cry_8_RNO_cZ(.I0(ZFF_X0_11_rep1),.I1(ZFF_X0[3:3]),.I2(ZFF_X0[13:13]),.O(un6_0_8_cry_8_RNO));
defparam un6_0_8_cry_8_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_8_cry_9_RNO_cZ(.I0(ZFF_X0_12_rep1),.I1(ZFF_X0[4:4]),.I2(ZFF_X0_14_rep1),.O(un6_0_8_cry_9_RNO));
defparam un6_0_8_cry_9_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_8_cry_10_RNO_cZ(.I0(ZFF_X0_fast[0:0]),.I1(ZFF_X0_15_rep1),.I2(ZFF_X0[5:5]),.O(un6_0_8_cry_10_RNO));
defparam un6_0_8_cry_10_RNO_cZ.INIT=8'h69;
  LUT3 un6_0_8_cry_13_RNO_cZ(.I0(ZFF_X0_fast[3:3]),.I1(ZFF_X0_fast[8:8]),.I2(ZFF_X0_fast[16:16]),.O(un6_0_8_cry_13_RNO));
defparam un6_0_8_cry_13_RNO_cZ.INIT=8'h69;
  LUT5 desc490(.I0(ZFF_X0_fast[3:3]),.I1(ZFF_X0_4_rep1),.I2(ZFF_X0_fast[9:9]),.I3(ZFF_X0_fast[8:8]),.I4(ZFF_X0_fast[16:16]),.O(un6_0_8_axb_14));
defparam desc490.INIT=32'h693CC369;
  LUT3 un6_0_8_cry_14_RNO_cZ(.I0(ZFF_X0_fast[3:3]),.I1(ZFF_X0_fast[8:8]),.I2(ZFF_X0_fast[16:16]),.O(un6_0_8_cry_14_RNO));
defparam un6_0_8_cry_14_RNO_cZ.INIT=8'hB2;
  LUT5 ZFF_X0_4_rep1_RNI6UT01(.I0(ZFF_X0_4_rep1),.I1(ZFF_X0_10_rep1),.I2(ZFF_X0_fast[9:9]),.I3(ZFF_X0_fast[5:5]),.I4(ZFF_X0_fast[16:16]),.O(un6_0_8_axb_15));
defparam ZFF_X0_4_rep1_RNI6UT01.INIT=32'h39C6C639;
  LUT2 un6_0_8_cry_15_RNO(.I0(ZFF_X0_4_rep1),.I1(ZFF_X0_fast[9:9]),.O(un6_0_6_1_scalar));
defparam un6_0_8_cry_15_RNO.INIT=4'h2;
  LUT3 un6_0_8_cry_16_RNO_cZ(.I0(ZFF_X0_10_rep1),.I1(ZFF_X0_fast[5:5]),.I2(ZFF_X0_fast[16:16]),.O(un6_0_8_cry_16_RNO));
defparam un6_0_8_cry_16_RNO_cZ.INIT=8'hD4;
  LUT5 ZFF_X0_11_rep1_RNIN8H21(.I0(ZFF_X0_11_rep1),.I1(ZFF_X0_6_rep1),.I2(ZFF_X0_7_rep1),.I3(ZFF_X0_12_rep1),.I4(ZFF_X0_fast[16:16]),.O(un6_0_8_axb_17));
defparam ZFF_X0_11_rep1_RNIN8H21.INIT=32'h4BB4B44B;
  LUT2 un6_0_8_cry_17_RNO_cZ(.I0(ZFF_X0_11_rep1),.I1(ZFF_X0_6_rep1),.O(un6_0_8_cry_17_RNO));
defparam un6_0_8_cry_17_RNO_cZ.INIT=4'h4;
  LUT5 desc491(.I0(ZFF_X0_fast[13:13]),.I1(ZFF_X0_7_rep1),.I2(ZFF_X0_12_rep1),.I3(ZFF_X0_fast[8:8]),.I4(ZFF_X0_fast[16:16]),.O(un6_0_8_axb_18));
defparam desc491.INIT=32'h659AA659;
  LUT3 un6_0_8_cry_18_RNO_cZ(.I0(ZFF_X0_7_rep1),.I1(ZFF_X0_12_rep1),.I2(ZFF_X0_fast[16:16]),.O(un6_0_8_cry_18_RNO));
defparam un6_0_8_cry_18_RNO_cZ.INIT=8'hB2;
  LUT5 desc492(.I0(ZFF_X0_fast[13:13]),.I1(ZFF_X0_14_rep1),.I2(ZFF_X0_fast[8:8]),.I3(ZFF_X0_fast[16:16]),.I4(ZFF_X0[9:9]),.O(un6_0_8_axb_19));
defparam desc492.INIT=32'h639C9C63;
  LUT2 un6_0_8_cry_19_RNO_cZ(.I0(ZFF_X0_fast[13:13]),.I1(ZFF_X0_fast[8:8]),.O(un6_0_8_cry_19_RNO));
defparam un6_0_8_cry_19_RNO_cZ.INIT=4'h4;
  LUT3 un6_0_8_cry_20_RNO_cZ(.I0(ZFF_X0_10_rep1),.I1(ZFF_X0_15_rep1),.I2(ZFF_X0_fast[16:16]),.O(un6_0_8_cry_20_RNO));
defparam un6_0_8_cry_20_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_8_cry_3_RNO_cZ(.I0(ZFF_X2_fast[6:6]),.I1(ZFF_X2_fast[8:8]),.I2(ZFF_X2_fast[5:5]),.O(un8_0_8_cry_3_RNO));
defparam un8_0_8_cry_3_RNO_cZ.INIT=8'h96;
  LUT3 un8_0_8_cry_4_RNO_cZ(.I0(ZFF_X2_fast[6:6]),.I1(ZFF_X2_fast[7:7]),.I2(ZFF_X2_fast[9:9]),.O(un8_0_8_cry_4_RNO));
defparam un8_0_8_cry_4_RNO_cZ.INIT=8'h96;
  LUT3 un8_0_8_cry_6_RNO_cZ(.I0(ZFF_X2_fast[1:1]),.I1(ZFF_X2_fast[11:11]),.I2(ZFF_X2_fast[9:9]),.O(un8_0_8_cry_6_RNO));
defparam un8_0_8_cry_6_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_8_cry_7_RNO_cZ(.I0(ZFF_X2[2:2]),.I1(ZFF_X2_10_rep1),.I2(ZFF_X2[12:12]),.O(un8_0_8_cry_7_RNO));
defparam un8_0_8_cry_7_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_8_cry_8_RNO_cZ(.I0(ZFF_X2_3_rep1),.I1(ZFF_X2[13:13]),.I2(ZFF_X2[11:11]),.O(un8_0_8_cry_8_RNO));
defparam un8_0_8_cry_8_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_8_cry_9_RNO_cZ(.I0(ZFF_X2_14_rep1),.I1(ZFF_X2[4:4]),.I2(ZFF_X2[12:12]),.O(un8_0_8_cry_9_RNO));
defparam un8_0_8_cry_9_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_8_cry_10_RNO_cZ(.I0(ZFF_X2_15_rep1),.I1(ZFF_X2[0:0]),.I2(ZFF_X2[5:5]),.O(un8_0_8_cry_10_RNO));
defparam un8_0_8_cry_10_RNO_cZ.INIT=8'h69;
  LUT3 un8_0_8_cry_13_RNO_cZ(.I0(ZFF_X2_fast[3:3]),.I1(ZFF_X2_fast[8:8]),.I2(ZFF_X2_fast[16:16]),.O(un8_0_8_cry_13_RNO));
defparam un8_0_8_cry_13_RNO_cZ.INIT=8'h69;
  LUT5 desc493(.I0(ZFF_X2_fast[3:3]),.I1(ZFF_X2_fast[8:8]),.I2(ZFF_X2_fast[4:4]),.I3(ZFF_X2_fast[9:9]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_8_axb_14));
defparam desc493.INIT=32'h4BB4D22D;
  LUT3 un8_0_8_cry_14_RNO_cZ(.I0(ZFF_X2_fast[3:3]),.I1(ZFF_X2_fast[8:8]),.I2(ZFF_X2_fast[16:16]),.O(un8_0_8_cry_14_RNO));
defparam un8_0_8_cry_14_RNO_cZ.INIT=8'hB2;
  LUT5 desc494(.I0(ZFF_X2_10_rep1),.I1(ZFF_X2_fast[4:4]),.I2(ZFF_X2_fast[9:9]),.I3(ZFF_X2_fast[5:5]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_8_axb_15));
defparam desc494.INIT=32'h59A6A659;
  LUT2 un8_0_8_cry_15_RNO(.I0(ZFF_X2_fast[4:4]),.I1(ZFF_X2_fast[9:9]),.O(un8_0_6_1_scalar));
defparam un8_0_8_cry_15_RNO.INIT=4'h2;
  LUT3 un8_0_8_cry_16_RNO_cZ(.I0(ZFF_X2_10_rep1),.I1(ZFF_X2_fast[5:5]),.I2(ZFF_X2_fast[16:16]),.O(un8_0_8_cry_16_RNO));
defparam un8_0_8_cry_16_RNO_cZ.INIT=8'hD4;
  LUT5 ZFF_X2_6_rep1_RNI1S1N(.I0(ZFF_X2_6_rep1),.I1(ZFF_X2_fast[11:11]),.I2(ZFF_X2_fast[12:12]),.I3(ZFF_X2[7:7]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_8_axb_17));
defparam ZFF_X2_6_rep1_RNI1S1N.INIT=32'h2DD2D22D;
  LUT2 un8_0_8_cry_17_RNO_cZ(.I0(ZFF_X2_6_rep1),.I1(ZFF_X2_fast[11:11]),.O(un8_0_8_cry_17_RNO));
defparam un8_0_8_cry_17_RNO_cZ.INIT=4'h2;
  LUT5 desc495(.I0(ZFF_X2_fast[13:13]),.I1(ZFF_X2_fast[12:12]),.I2(ZFF_X2[7:7]),.I3(ZFF_X2[8:8]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_8_axb_18));
defparam desc495.INIT=32'h59A69A65;
  LUT3 un8_0_8_cry_18_RNO_cZ(.I0(ZFF_X2_fast[12:12]),.I1(ZFF_X2[7:7]),.I2(ZFF_X2_fast[16:16]),.O(un8_0_8_cry_18_RNO));
defparam un8_0_8_cry_18_RNO_cZ.INIT=8'hD4;
  LUT5 desc496(.I0(ZFF_X2_fast[13:13]),.I1(ZFF_X2_14_rep1),.I2(ZFF_X2[9:9]),.I3(ZFF_X2[8:8]),.I4(ZFF_X2_fast[16:16]),.O(un8_0_8_axb_19));
defparam desc496.INIT=32'h693C96C3;
  LUT2 un8_0_8_cry_19_RNO_cZ(.I0(ZFF_X2_fast[13:13]),.I1(ZFF_X2[8:8]),.O(un8_0_8_cry_19_RNO));
defparam un8_0_8_cry_19_RNO_cZ.INIT=4'h4;
  LUT3 un8_0_8_cry_20_RNO_cZ(.I0(ZFF_X2_15_rep1),.I1(ZFF_X2_10_rep1),.I2(ZFF_X2_fast[16:16]),.O(un8_0_8_cry_20_RNO));
defparam un8_0_8_cry_20_RNO_cZ.INIT=8'h69;
  LUT2 un10_8_cry_11_RNO_cZ(.I0(ZFF_Y2[0:0]),.I1(ZFF_Y2[2:2]),.O(un10_8_cry_11_RNO));
defparam un10_8_cry_11_RNO_cZ.INIT=4'h8;
  LUT3 Y_out_double_2_6_0_s_0_RNIQS6I(.I0(pgZFF_X0[0:0]),.I1(pgZFF_X2[0:0]),.I2(Y_out_double_2_6[0:0]),.O(Y_out_double_2[0:0]));
defparam Y_out_double_2_6_0_s_0_RNIQS6I.INIT=8'h96;
  LUT2 desc497(.I0(pgZFF_X0[0:0]),.I1(pgZFF_X2[0:0]),.O(Y_out_double_2_4[0:0]));
defparam desc497.INIT=4'h6;
  XORCY Y_out_double_2_4_s_17(.LI(Y_out_double_2_4_axb_17),.CI(Y_out_double_2_4_cry_16),.O(Y_out_double_2_4[17:17]));
  XORCY Y_out_double_2_4_s_16(.LI(Y_out_double_2_4_axb_16),.CI(Y_out_double_2_4_cry_15),.O(Y_out_double_2_4[16:16]));
  MUXCY_L Y_out_double_2_4_cry_16_cZ(.DI(Y_out_double_2_7[17:17]),.CI(Y_out_double_2_4_cry_15),.S(Y_out_double_2_4_axb_16),.LO(Y_out_double_2_4_cry_16));
  XORCY Y_out_double_2_4_s_15(.LI(Y_out_double_2_4_axb_15),.CI(Y_out_double_2_4_cry_14),.O(Y_out_double_2_4[15:15]));
  MUXCY_L Y_out_double_2_4_cry_15_cZ(.DI(Y_out_double_2_7[15:15]),.CI(Y_out_double_2_4_cry_14),.S(Y_out_double_2_4_axb_15),.LO(Y_out_double_2_4_cry_15));
  XORCY Y_out_double_2_4_s_14(.LI(Y_out_double_2_4_axb_14),.CI(Y_out_double_2_4_cry_13),.O(Y_out_double_2_4[14:14]));
  MUXCY_L Y_out_double_2_4_cry_14_cZ(.DI(Y_out_double_2_7[14:14]),.CI(Y_out_double_2_4_cry_13),.S(Y_out_double_2_4_axb_14),.LO(Y_out_double_2_4_cry_14));
  XORCY Y_out_double_2_4_s_13(.LI(Y_out_double_2_4_axb_13),.CI(Y_out_double_2_4_cry_12),.O(Y_out_double_2_4[13:13]));
  MUXCY_L Y_out_double_2_4_cry_13_cZ(.DI(Y_out_double_2_7[13:13]),.CI(Y_out_double_2_4_cry_12),.S(Y_out_double_2_4_axb_13),.LO(Y_out_double_2_4_cry_13));
  XORCY Y_out_double_2_4_s_12(.LI(Y_out_double_2_4_axb_12),.CI(Y_out_double_2_4_cry_11),.O(Y_out_double_2_4[12:12]));
  MUXCY_L Y_out_double_2_4_cry_12_cZ(.DI(Y_out_double_2_7[12:12]),.CI(Y_out_double_2_4_cry_11),.S(Y_out_double_2_4_axb_12),.LO(Y_out_double_2_4_cry_12));
  XORCY Y_out_double_2_4_s_11(.LI(Y_out_double_2_4_axb_11),.CI(Y_out_double_2_4_cry_10),.O(Y_out_double_2_4[11:11]));
  MUXCY_L Y_out_double_2_4_cry_11_cZ(.DI(Y_out_double_2_7[11:11]),.CI(Y_out_double_2_4_cry_10),.S(Y_out_double_2_4_axb_11),.LO(Y_out_double_2_4_cry_11));
  XORCY Y_out_double_2_4_s_10(.LI(Y_out_double_2_4_axb_10),.CI(Y_out_double_2_4_cry_9),.O(Y_out_double_2_4[10:10]));
  MUXCY_L Y_out_double_2_4_cry_10_cZ(.DI(Y_out_double_2_7[10:10]),.CI(Y_out_double_2_4_cry_9),.S(Y_out_double_2_4_axb_10),.LO(Y_out_double_2_4_cry_10));
  XORCY Y_out_double_2_4_s_9(.LI(Y_out_double_2_4_axb_9),.CI(Y_out_double_2_4_cry_8),.O(Y_out_double_2_4[9:9]));
  MUXCY_L Y_out_double_2_4_cry_9_cZ(.DI(Y_out_double_2_7[9:9]),.CI(Y_out_double_2_4_cry_8),.S(Y_out_double_2_4_axb_9),.LO(Y_out_double_2_4_cry_9));
  XORCY Y_out_double_2_4_s_8(.LI(Y_out_double_2_4_axb_8),.CI(Y_out_double_2_4_cry_7),.O(Y_out_double_2_4[8:8]));
  MUXCY_L Y_out_double_2_4_cry_8_cZ(.DI(Y_out_double_2_7[8:8]),.CI(Y_out_double_2_4_cry_7),.S(Y_out_double_2_4_axb_8),.LO(Y_out_double_2_4_cry_8));
  XORCY Y_out_double_2_4_s_7(.LI(Y_out_double_2_4_axb_7),.CI(Y_out_double_2_4_cry_6),.O(Y_out_double_2_4[7:7]));
  MUXCY_L Y_out_double_2_4_cry_7_cZ(.DI(Y_out_double_2_7[7:7]),.CI(Y_out_double_2_4_cry_6),.S(Y_out_double_2_4_axb_7),.LO(Y_out_double_2_4_cry_7));
  XORCY Y_out_double_2_4_s_6(.LI(Y_out_double_2_4_axb_6),.CI(Y_out_double_2_4_cry_5),.O(Y_out_double_2_4[6:6]));
  MUXCY_L Y_out_double_2_4_cry_6_cZ(.DI(Y_out_double_2_7[6:6]),.CI(Y_out_double_2_4_cry_5),.S(Y_out_double_2_4_axb_6),.LO(Y_out_double_2_4_cry_6));
  XORCY Y_out_double_2_4_s_5(.LI(Y_out_double_2_4_axb_5),.CI(Y_out_double_2_4_cry_4),.O(Y_out_double_2_4[5:5]));
  MUXCY_L Y_out_double_2_4_cry_5_cZ(.DI(Y_out_double_2_7[5:5]),.CI(Y_out_double_2_4_cry_4),.S(Y_out_double_2_4_axb_5),.LO(Y_out_double_2_4_cry_5));
  XORCY Y_out_double_2_4_s_4(.LI(Y_out_double_2_4_axb_4),.CI(Y_out_double_2_4_cry_3),.O(Y_out_double_2_4[4:4]));
  MUXCY_L Y_out_double_2_4_cry_4_cZ(.DI(Y_out_double_2_7[4:4]),.CI(Y_out_double_2_4_cry_3),.S(Y_out_double_2_4_axb_4),.LO(Y_out_double_2_4_cry_4));
  XORCY Y_out_double_2_4_s_3(.LI(Y_out_double_2_4_axb_3),.CI(Y_out_double_2_4_cry_2),.O(Y_out_double_2_4[3:3]));
  MUXCY_L Y_out_double_2_4_cry_3_cZ(.DI(Y_out_double_2_7[3:3]),.CI(Y_out_double_2_4_cry_2),.S(Y_out_double_2_4_axb_3),.LO(Y_out_double_2_4_cry_3));
  XORCY Y_out_double_2_4_s_2(.LI(Y_out_double_2_4_axb_2),.CI(Y_out_double_2_4_cry_1),.O(Y_out_double_2_4[2:2]));
  MUXCY_L Y_out_double_2_4_cry_2_cZ(.DI(Y_out_double_2_7[2:2]),.CI(Y_out_double_2_4_cry_1),.S(Y_out_double_2_4_axb_2),.LO(Y_out_double_2_4_cry_2));
  XORCY Y_out_double_2_4_s_1(.LI(Y_out_double_2_4_axb_1),.CI(Y_out_double_2_4_cry_0),.O(Y_out_double_2_4[1:1]));
  MUXCY_L Y_out_double_2_4_cry_1_cZ(.DI(pgZFF_X2[1:1]),.CI(Y_out_double_2_4_cry_0),.S(Y_out_double_2_4_axb_1),.LO(Y_out_double_2_4_cry_1));
  MUXCY_L Y_out_double_2_4_cry_0_cZ(.DI(pgZFF_X2[0:0]),.CI(GND),.S(Y_out_double_2_4[0:0]),.LO(Y_out_double_2_4_cry_0));
  XORCY un9_11_s_24(.LI(un9_11_axb_24),.CI(un9_11_cry_23),.O(un9_11[45:45]));
  MUXCY un9_11_cry_24(.DI(GND),.CI(un9_11_cry_23),.S(un9_11_axb_24),.O(un9_11_0[46:46]));
  XORCY un9_11_s_23(.LI(un9_11_axb_23),.CI(un9_11_cry_22),.O(un9_11[44:44]));
  MUXCY_L un9_11_cry_23_cZ(.DI(GND),.CI(un9_11_cry_22),.S(un9_11_axb_23),.LO(un9_11_cry_23));
  XORCY un9_11_s_22(.LI(un9_11_axb_22),.CI(un9_11_cry_21),.O(un9_11[43:43]));
  MUXCY_L un9_11_cry_22_cZ(.DI(ZFF_Y1_16_rep1),.CI(un9_11_cry_21),.S(un9_11_axb_22),.LO(un9_11_cry_22));
  XORCY un9_11_s_21(.LI(un9_11_axb_21),.CI(un9_11_cry_20),.O(un9_11[42:42]));
  MUXCY_L un9_11_cry_21_cZ(.DI(ZFF_Y1_15_rep1),.CI(un9_11_cry_20),.S(un9_11_axb_21),.LO(un9_11_cry_21));
  XORCY un9_11_s_20(.LI(un9_11_axb_20),.CI(un9_11_cry_19),.O(un9_11[41:41]));
  MUXCY_L un9_11_cry_20_cZ(.DI(un9_11_26_rep1),.CI(un9_11_cry_19),.S(un9_11_axb_20),.LO(un9_11_cry_20));
  XORCY un9_11_s_19(.LI(un9_11_axb_19),.CI(un9_11_cry_18),.O(un9_11[40:40]));
  MUXCY_L un9_11_cry_19_cZ(.DI(un9_11_25_rep1),.CI(un9_11_cry_18),.S(un9_11_axb_19),.LO(un9_11_cry_19));
  XORCY un9_11_s_18(.LI(un9_11_axb_18),.CI(un9_11_cry_17),.O(un9_11[39:39]));
  MUXCY_L un9_11_cry_18_cZ(.DI(un9_11_fast[24:24]),.CI(un9_11_cry_17),.S(un9_11_axb_18),.LO(un9_11_cry_18));
  XORCY un9_11_s_17(.LI(un9_11_axb_17),.CI(un9_11_cry_16),.O(un9_11[38:38]));
  MUXCY_L un9_11_cry_17_cZ(.DI(un9_11_fast[23:23]),.CI(un9_11_cry_16),.S(un9_11_axb_17),.LO(un9_11_cry_17));
  XORCY un9_11_s_16(.LI(un9_11_axb_16),.CI(un9_11_cry_15),.O(un9_11[37:37]));
  MUXCY_L un9_11_cry_16_cZ(.DI(un9_11_fast[22:22]),.CI(un9_11_cry_15),.S(un9_11_axb_16),.LO(un9_11_cry_16));
  XORCY un9_11_s_15(.LI(un9_11_axb_15),.CI(un9_11_cry_14),.O(un9_11[36:36]));
  MUXCY_L un9_11_cry_15_cZ(.DI(ZFF_Y1_fast[9:9]),.CI(un9_11_cry_14),.S(un9_11_axb_15),.LO(un9_11_cry_15));
  XORCY un9_11_s_14(.LI(un9_11_axb_14),.CI(un9_11_cry_13),.O(un9_11[35:35]));
  MUXCY_L un9_11_cry_14_cZ(.DI(ZFF_Y1_fast[8:8]),.CI(un9_11_cry_13),.S(un9_11_axb_14),.LO(un9_11_cry_14));
  XORCY un9_11_s_13(.LI(un9_11_axb_13),.CI(un9_11_cry_12),.O(un9_11[34:34]));
  MUXCY_L un9_11_cry_13_cZ(.DI(ZFF_Y1_fast[7:7]),.CI(un9_11_cry_12),.S(un9_11_axb_13),.LO(un9_11_cry_13));
  XORCY un9_11_s_12(.LI(un9_11_axb_12),.CI(un9_11_cry_11),.O(un9_11[33:33]));
  MUXCY_L un9_11_cry_12_cZ(.DI(ZFF_Y1_fast[6:6]),.CI(un9_11_cry_11),.S(un9_11_axb_12),.LO(un9_11_cry_12));
  XORCY un9_11_s_11(.LI(un9_11_axb_11),.CI(un9_11_cry_10),.O(un9_11[32:32]));
  MUXCY_L un9_11_cry_11_cZ(.DI(ZFF_Y1_fast[5:5]),.CI(un9_11_cry_10),.S(un9_11_axb_11),.LO(un9_11_cry_11));
  XORCY un9_11_s_10(.LI(un9_11_axb_10),.CI(un9_11_cry_9),.O(un9_11[31:31]));
  MUXCY_L un9_11_cry_10_cZ(.DI(ZFF_Y1_fast[4:4]),.CI(un9_11_cry_9),.S(un9_11_axb_10),.LO(un9_11_cry_10));
  XORCY un9_11_s_9(.LI(un9_11_axb_9),.CI(un9_11_cry_8),.O(un9_11[30:30]));
  MUXCY_L un9_11_cry_9_cZ(.DI(ZFF_Y1_fast[3:3]),.CI(un9_11_cry_8),.S(un9_11_axb_9),.LO(un9_11_cry_9));
  XORCY un9_11_s_8(.LI(un9_11_axb_8),.CI(un9_11_cry_7),.O(un9_11[29:29]));
  MUXCY_L un9_11_cry_8_cZ(.DI(un9_8_fast[7:7]),.CI(un9_11_cry_7),.S(un9_11_axb_8),.LO(un9_11_cry_8));
  XORCY un9_11_s_7(.LI(un9_11_axb_7),.CI(un9_11_cry_6),.O(un9_11[28:28]));
  MUXCY_L un9_11_cry_7_cZ(.DI(ZFF_Y1_fast[16:16]),.CI(un9_11_cry_6),.S(un9_11_axb_7),.LO(un9_11_cry_7));
  MUXCY_L un9_11_cry_6_cZ(.DI(ZFF_Y1_fast[15:15]),.CI(GND),.S(un9_11_cry_6_RNO),.LO(un9_11_cry_6));
  XORCY un8_0_9_s_26(.LI(un8_0_9_axb_26),.CI(un8_0_9_cry_25),.O(un8_0_9[41:41]));
  MUXCY un8_0_9_cry_26(.DI(GND),.CI(un8_0_9_cry_25),.S(un8_0_9_axb_26),.O(un8_0_9_0[42:42]));
  XORCY un8_0_9_s_25(.LI(un8_0_9_axb_25),.CI(un8_0_9_cry_24),.O(un8_0_9[40:40]));
  MUXCY_L un8_0_9_cry_25_cZ(.DI(GND),.CI(un8_0_9_cry_24),.S(un8_0_9_axb_25),.LO(un8_0_9_cry_25));
  XORCY un8_0_9_s_24(.LI(un8_0_9_axb_24),.CI(un8_0_9_cry_23),.O(un8_0_9[39:39]));
  MUXCY_L un8_0_9_cry_24_cZ(.DI(GND),.CI(un8_0_9_cry_23),.S(un8_0_9_axb_24),.LO(un8_0_9_cry_24));
  XORCY un8_0_9_s_23(.LI(un8_0_9_axb_23),.CI(un8_0_9_cry_22),.O(un8_0_9[38:38]));
  MUXCY_L un8_0_9_cry_23_cZ(.DI(ZFF_X2[12:12]),.CI(un8_0_9_cry_22),.S(un8_0_9_axb_23),.LO(un8_0_9_cry_23));
  XORCY un8_0_9_s_22(.LI(un8_0_9_axb_22),.CI(un8_0_9_cry_21),.O(un8_0_9[37:37]));
  MUXCY_L un8_0_9_cry_22_cZ(.DI(ZFF_X2[11:11]),.CI(un8_0_9_cry_21),.S(un8_0_9_axb_22),.LO(un8_0_9_cry_22));
  XORCY un8_0_9_s_21(.LI(un8_0_9_axb_21),.CI(un8_0_9_cry_20),.O(un8_0_9[36:36]));
  MUXCY_L un8_0_9_cry_21_cZ(.DI(ZFF_X2[10:10]),.CI(un8_0_9_cry_20),.S(un8_0_9_axb_21),.LO(un8_0_9_cry_21));
  XORCY un8_0_9_s_20(.LI(un8_0_9_axb_20),.CI(un8_0_9_cry_19),.O(un8_0_9[35:35]));
  MUXCY_L un8_0_9_cry_20_cZ(.DI(ZFF_X2[9:9]),.CI(un8_0_9_cry_19),.S(un8_0_9_axb_20),.LO(un8_0_9_cry_20));
  XORCY un8_0_9_s_19(.LI(un8_0_9_axb_19),.CI(un8_0_9_cry_18),.O(un8_0_9[34:34]));
  MUXCY_L un8_0_9_cry_19_cZ(.DI(ZFF_X2[8:8]),.CI(un8_0_9_cry_18),.S(un8_0_9_axb_19),.LO(un8_0_9_cry_19));
  XORCY un8_0_9_s_18(.LI(un8_0_9_axb_18),.CI(un8_0_9_cry_17),.O(un8_0_9[33:33]));
  MUXCY_L un8_0_9_cry_18_cZ(.DI(ZFF_X2[7:7]),.CI(un8_0_9_cry_17),.S(un8_0_9_axb_18),.LO(un8_0_9_cry_18));
  XORCY un8_0_9_s_17(.LI(un8_0_9_axb_17),.CI(un8_0_9_cry_16),.O(un8_0_9[32:32]));
  MUXCY_L un8_0_9_cry_17_cZ(.DI(ZFF_X2[6:6]),.CI(un8_0_9_cry_16),.S(un8_0_9_axb_17),.LO(un8_0_9_cry_17));
  XORCY un8_0_9_s_16(.LI(un8_0_9_axb_16),.CI(un8_0_9_cry_15),.O(un8_0_9[31:31]));
  MUXCY_L un8_0_9_cry_16_cZ(.DI(ZFF_X2[5:5]),.CI(un8_0_9_cry_15),.S(un8_0_9_axb_16),.LO(un8_0_9_cry_16));
  XORCY un8_0_9_s_15(.LI(un8_0_9_axb_15),.CI(un8_0_9_cry_14),.O(un8_0_9[30:30]));
  MUXCY_L un8_0_9_cry_15_cZ(.DI(ZFF_X2[4:4]),.CI(un8_0_9_cry_14),.S(un8_0_9_axb_15),.LO(un8_0_9_cry_15));
  XORCY un8_0_9_s_14(.LI(un8_0_9_axb_14),.CI(un8_0_9_cry_13),.O(un8_0_9[29:29]));
  MUXCY_L un8_0_9_cry_14_cZ(.DI(ZFF_X2[3:3]),.CI(un8_0_9_cry_13),.S(un8_0_9_axb_14),.LO(un8_0_9_cry_14));
  XORCY un8_0_9_s_13(.LI(un8_0_9_axb_13),.CI(un8_0_9_cry_12),.O(un8_0_9[28:28]));
  MUXCY_L un8_0_9_cry_13_cZ(.DI(ZFF_X2[2:2]),.CI(un8_0_9_cry_12),.S(un8_0_9_axb_13),.LO(un8_0_9_cry_13));
  XORCY un8_0_9_s_12(.LI(un8_0_9_axb_12),.CI(un8_0_9_cry_11),.O(un8_0_9[27:27]));
  MUXCY_L un8_0_9_cry_12_cZ(.DI(ZFF_X2[1:1]),.CI(un8_0_9_cry_11),.S(un8_0_9_axb_12),.LO(un8_0_9_cry_12));
  XORCY un8_0_9_s_11(.LI(un8_0_9_axb_11),.CI(un8_0_9_cry_10),.O(un8_0_9[26:26]));
  MUXCY_L un8_0_9_cry_11_cZ(.DI(ZFF_X2[0:0]),.CI(un8_0_9_cry_10),.S(un8_0_9_axb_11),.LO(un8_0_9_cry_11));
  XORCY un8_0_9_s_10(.LI(un8_0_9_axb_10),.CI(un8_0_9_cry_9),.O(un8_0_9[25:25]));
  MUXCY_L un8_0_9_cry_10_cZ(.DI(GND),.CI(un8_0_9_cry_9),.S(un8_0_9_axb_10),.LO(un8_0_9_cry_10));
  XORCY un8_0_9_s_9(.LI(un8_0_9_axb_9),.CI(un8_0_9_cry_8),.O(un8_0_9[24:24]));
  MUXCY_L un8_0_9_cry_9_cZ(.DI(GND),.CI(un8_0_9_cry_8),.S(un8_0_9_axb_9),.LO(un8_0_9_cry_9));
  XORCY un8_0_9_s_8(.LI(un8_0_9_axb_8),.CI(un8_0_9_cry_7),.O(un8_0_9[23:23]));
  MUXCY_L un8_0_9_cry_8_cZ(.DI(GND),.CI(un8_0_9_cry_7),.S(un8_0_9_axb_8),.LO(un8_0_9_cry_8));
  XORCY un8_0_9_s_7(.LI(un8_0_9_axb_7),.CI(un8_0_9_cry_6),.O(un8_0_9[22:22]));
  MUXCY_L un8_0_9_cry_7_cZ(.DI(GND),.CI(un8_0_9_cry_6),.S(un8_0_9_axb_7),.LO(un8_0_9_cry_7));
  XORCY un8_0_9_s_6(.LI(un8_0_9_axb_6),.CI(un8_0_9_cry_5),.O(un8_0_9[21:21]));
  MUXCY_L un8_0_9_cry_6_cZ(.DI(GND),.CI(un8_0_9_cry_5),.S(un8_0_9_axb_6),.LO(un8_0_9_cry_6));
  XORCY un8_0_9_s_5(.LI(un8_0_9_axb_5),.CI(un8_0_9_cry_4),.O(un8_0_9[20:20]));
  MUXCY_L un8_0_9_cry_5_cZ(.DI(ZFF_X2[12:12]),.CI(un8_0_9_cry_4),.S(un8_0_9_axb_5),.LO(un8_0_9_cry_5));
  XORCY un8_0_9_s_4(.LI(un8_0_9_axb_4),.CI(un8_0_9_cry_3),.O(un8_0_9[19:19]));
  MUXCY_L un8_0_9_cry_4_cZ(.DI(GND),.CI(un8_0_9_cry_3),.S(un8_0_9_axb_4),.LO(un8_0_9_cry_4));
  XORCY un8_0_9_s_3(.LI(un8_0_9_axb_3),.CI(un8_0_9_cry_2),.O(un8_0_9[18:18]));
  MUXCY_L un8_0_9_cry_3_cZ(.DI(GND),.CI(un8_0_9_cry_2),.S(un8_0_9_axb_3),.LO(un8_0_9_cry_3));
  XORCY un8_0_9_s_2(.LI(un8_0_9_axb_2),.CI(un8_0_9_cry_1),.O(un8_0_9[17:17]));
  MUXCY_L un8_0_9_cry_2_cZ(.DI(GND),.CI(un8_0_9_cry_1),.S(un8_0_9_axb_2),.LO(un8_0_9_cry_2));
  XORCY un8_0_9_s_1(.LI(un8_0_9_axb_1),.CI(un8_0_9_cry_0),.O(un8_0_9[16:16]));
  MUXCY_L un8_0_9_cry_1_cZ(.DI(GND),.CI(un8_0_9_cry_0),.S(un8_0_9_axb_1),.LO(un8_0_9_cry_1));
  MUXCY_L un8_0_9_cry_0_cZ(.DI(ZFF_X2_fast[7:7]),.CI(GND),.S(un8_0_9[15:15]),.LO(un8_0_9_cry_0));
  XORCY un6_0_9_s_26(.LI(un6_0_9_axb_26),.CI(un6_0_9_cry_25),.O(un6_0_9[41:41]));
  MUXCY un6_0_9_cry_26(.DI(GND),.CI(un6_0_9_cry_25),.S(un6_0_9_axb_26),.O(un6_0_9_0[42:42]));
  XORCY un6_0_9_s_25(.LI(un6_0_9_axb_25),.CI(un6_0_9_cry_24),.O(un6_0_9[40:40]));
  MUXCY_L un6_0_9_cry_25_cZ(.DI(GND),.CI(un6_0_9_cry_24),.S(un6_0_9_axb_25),.LO(un6_0_9_cry_25));
  XORCY un6_0_9_s_24(.LI(un6_0_9_axb_24),.CI(un6_0_9_cry_23),.O(un6_0_9[39:39]));
  MUXCY_L un6_0_9_cry_24_cZ(.DI(GND),.CI(un6_0_9_cry_23),.S(un6_0_9_axb_24),.LO(un6_0_9_cry_24));
  XORCY un6_0_9_s_23(.LI(un6_0_9_axb_23),.CI(un6_0_9_cry_22),.O(un6_0_9[38:38]));
  MUXCY_L un6_0_9_cry_23_cZ(.DI(ZFF_X0[12:12]),.CI(un6_0_9_cry_22),.S(un6_0_9_axb_23),.LO(un6_0_9_cry_23));
  XORCY un6_0_9_s_22(.LI(un6_0_9_axb_22),.CI(un6_0_9_cry_21),.O(un6_0_9[37:37]));
  MUXCY_L un6_0_9_cry_22_cZ(.DI(ZFF_X0[11:11]),.CI(un6_0_9_cry_21),.S(un6_0_9_axb_22),.LO(un6_0_9_cry_22));
  XORCY un6_0_9_s_21(.LI(un6_0_9_axb_21),.CI(un6_0_9_cry_20),.O(un6_0_9[36:36]));
  MUXCY_L un6_0_9_cry_21_cZ(.DI(ZFF_X0[10:10]),.CI(un6_0_9_cry_20),.S(un6_0_9_axb_21),.LO(un6_0_9_cry_21));
  XORCY un6_0_9_s_20(.LI(un6_0_9_axb_20),.CI(un6_0_9_cry_19),.O(un6_0_9[35:35]));
  MUXCY_L un6_0_9_cry_20_cZ(.DI(ZFF_X0[9:9]),.CI(un6_0_9_cry_19),.S(un6_0_9_axb_20),.LO(un6_0_9_cry_20));
  XORCY un6_0_9_s_19(.LI(un6_0_9_axb_19),.CI(un6_0_9_cry_18),.O(un6_0_9[34:34]));
  MUXCY_L un6_0_9_cry_19_cZ(.DI(ZFF_X0[8:8]),.CI(un6_0_9_cry_18),.S(un6_0_9_axb_19),.LO(un6_0_9_cry_19));
  XORCY un6_0_9_s_18(.LI(un6_0_9_axb_18),.CI(un6_0_9_cry_17),.O(un6_0_9[33:33]));
  MUXCY_L un6_0_9_cry_18_cZ(.DI(ZFF_X0[7:7]),.CI(un6_0_9_cry_17),.S(un6_0_9_axb_18),.LO(un6_0_9_cry_18));
  XORCY un6_0_9_s_17(.LI(un6_0_9_axb_17),.CI(un6_0_9_cry_16),.O(un6_0_9[32:32]));
  MUXCY_L un6_0_9_cry_17_cZ(.DI(ZFF_X0[6:6]),.CI(un6_0_9_cry_16),.S(un6_0_9_axb_17),.LO(un6_0_9_cry_17));
  XORCY un6_0_9_s_16(.LI(un6_0_9_axb_16),.CI(un6_0_9_cry_15),.O(un6_0_9[31:31]));
  MUXCY_L un6_0_9_cry_16_cZ(.DI(ZFF_X0[5:5]),.CI(un6_0_9_cry_15),.S(un6_0_9_axb_16),.LO(un6_0_9_cry_16));
  XORCY un6_0_9_s_15(.LI(un6_0_9_axb_15),.CI(un6_0_9_cry_14),.O(un6_0_9[30:30]));
  MUXCY_L un6_0_9_cry_15_cZ(.DI(ZFF_X0[4:4]),.CI(un6_0_9_cry_14),.S(un6_0_9_axb_15),.LO(un6_0_9_cry_15));
  XORCY un6_0_9_s_14(.LI(un6_0_9_axb_14),.CI(un6_0_9_cry_13),.O(un6_0_9[29:29]));
  MUXCY_L un6_0_9_cry_14_cZ(.DI(ZFF_X0[3:3]),.CI(un6_0_9_cry_13),.S(un6_0_9_axb_14),.LO(un6_0_9_cry_14));
  XORCY un6_0_9_s_13(.LI(un6_0_9_axb_13),.CI(un6_0_9_cry_12),.O(un6_0_9[28:28]));
  MUXCY_L un6_0_9_cry_13_cZ(.DI(ZFF_X0[2:2]),.CI(un6_0_9_cry_12),.S(un6_0_9_axb_13),.LO(un6_0_9_cry_13));
  XORCY un6_0_9_s_12(.LI(un6_0_9_axb_12),.CI(un6_0_9_cry_11),.O(un6_0_9[27:27]));
  MUXCY_L un6_0_9_cry_12_cZ(.DI(ZFF_X0[1:1]),.CI(un6_0_9_cry_11),.S(un6_0_9_axb_12),.LO(un6_0_9_cry_12));
  XORCY un6_0_9_s_11(.LI(un6_0_9_axb_11),.CI(un6_0_9_cry_10),.O(un6_0_9[26:26]));
  MUXCY_L un6_0_9_cry_11_cZ(.DI(ZFF_X0[0:0]),.CI(un6_0_9_cry_10),.S(un6_0_9_axb_11),.LO(un6_0_9_cry_11));
  XORCY un6_0_9_s_10(.LI(un6_0_9_axb_10),.CI(un6_0_9_cry_9),.O(un6_0_9[25:25]));
  MUXCY_L un6_0_9_cry_10_cZ(.DI(GND),.CI(un6_0_9_cry_9),.S(un6_0_9_axb_10),.LO(un6_0_9_cry_10));
  XORCY un6_0_9_s_9(.LI(un6_0_9_axb_9),.CI(un6_0_9_cry_8),.O(un6_0_9[24:24]));
  MUXCY_L un6_0_9_cry_9_cZ(.DI(GND),.CI(un6_0_9_cry_8),.S(un6_0_9_axb_9),.LO(un6_0_9_cry_9));
  XORCY un6_0_9_s_8(.LI(un6_0_9_axb_8),.CI(un6_0_9_cry_7),.O(un6_0_9[23:23]));
  MUXCY_L un6_0_9_cry_8_cZ(.DI(GND),.CI(un6_0_9_cry_7),.S(un6_0_9_axb_8),.LO(un6_0_9_cry_8));
  XORCY un6_0_9_s_7(.LI(un6_0_9_axb_7),.CI(un6_0_9_cry_6),.O(un6_0_9[22:22]));
  MUXCY_L un6_0_9_cry_7_cZ(.DI(GND),.CI(un6_0_9_cry_6),.S(un6_0_9_axb_7),.LO(un6_0_9_cry_7));
  XORCY un6_0_9_s_6(.LI(un6_0_9_axb_6),.CI(un6_0_9_cry_5),.O(un6_0_9[21:21]));
  MUXCY_L un6_0_9_cry_6_cZ(.DI(GND),.CI(un6_0_9_cry_5),.S(un6_0_9_axb_6),.LO(un6_0_9_cry_6));
  XORCY un6_0_9_s_5(.LI(un6_0_9_axb_5),.CI(un6_0_9_cry_4),.O(un6_0_9[20:20]));
  MUXCY_L un6_0_9_cry_5_cZ(.DI(ZFF_X0_12_rep1),.CI(un6_0_9_cry_4),.S(un6_0_9_axb_5),.LO(un6_0_9_cry_5));
  XORCY un6_0_9_s_4(.LI(un6_0_9_axb_4),.CI(un6_0_9_cry_3),.O(un6_0_9[19:19]));
  MUXCY_L un6_0_9_cry_4_cZ(.DI(GND),.CI(un6_0_9_cry_3),.S(un6_0_9_axb_4),.LO(un6_0_9_cry_4));
  XORCY un6_0_9_s_3(.LI(un6_0_9_axb_3),.CI(un6_0_9_cry_2),.O(un6_0_9[18:18]));
  MUXCY_L un6_0_9_cry_3_cZ(.DI(GND),.CI(un6_0_9_cry_2),.S(un6_0_9_axb_3),.LO(un6_0_9_cry_3));
  XORCY un6_0_9_s_2(.LI(un6_0_9_axb_2),.CI(un6_0_9_cry_1),.O(un6_0_9[17:17]));
  MUXCY_L un6_0_9_cry_2_cZ(.DI(GND),.CI(un6_0_9_cry_1),.S(un6_0_9_axb_2),.LO(un6_0_9_cry_2));
  XORCY un6_0_9_s_1(.LI(un6_0_9_axb_1),.CI(un6_0_9_cry_0),.O(un6_0_9[16:16]));
  MUXCY_L un6_0_9_cry_1_cZ(.DI(GND),.CI(un6_0_9_cry_0),.S(un6_0_9_axb_1),.LO(un6_0_9_cry_1));
  MUXCY_L un6_0_9_cry_0_cZ(.DI(ZFF_X0_fast[7:7]),.CI(GND),.S(un6_0_9[15:15]),.LO(un6_0_9_cry_0));
  XORCY Y_out_double_2_7_s_16(.LI(Y_out_double_2_7_axb_16),.CI(Y_out_double_2_7_cry_15),.O(Y_out_double_2_7[17:17]));
  XORCY Y_out_double_2_7_s_15(.LI(Y_out_double_2_7_axb_15),.CI(Y_out_double_2_7_cry_14),.O(Y_out_double_2_7[15:15]));
  MUXCY_L Y_out_double_2_7_cry_15_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_14),.S(Y_out_double_2_7_axb_15),.LO(Y_out_double_2_7_cry_15));
  XORCY Y_out_double_2_7_s_14(.LI(Y_out_double_2_7_axb_14),.CI(Y_out_double_2_7_cry_13),.O(Y_out_double_2_7[14:14]));
  MUXCY_L Y_out_double_2_7_cry_14_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_13),.S(Y_out_double_2_7_axb_14),.LO(Y_out_double_2_7_cry_14));
  XORCY Y_out_double_2_7_s_13(.LI(Y_out_double_2_7_axb_13),.CI(Y_out_double_2_7_cry_12),.O(Y_out_double_2_7[13:13]));
  MUXCY_L Y_out_double_2_7_cry_13_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_12),.S(Y_out_double_2_7_axb_13),.LO(Y_out_double_2_7_cry_13));
  XORCY Y_out_double_2_7_s_12(.LI(Y_out_double_2_7_axb_12),.CI(Y_out_double_2_7_cry_11),.O(Y_out_double_2_7[12:12]));
  MUXCY_L Y_out_double_2_7_cry_12_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_11),.S(Y_out_double_2_7_axb_12),.LO(Y_out_double_2_7_cry_12));
  XORCY Y_out_double_2_7_s_11(.LI(Y_out_double_2_7_axb_11),.CI(Y_out_double_2_7_cry_10),.O(Y_out_double_2_7[11:11]));
  MUXCY_L Y_out_double_2_7_cry_11_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_10),.S(Y_out_double_2_7_axb_11),.LO(Y_out_double_2_7_cry_11));
  XORCY Y_out_double_2_7_s_10(.LI(Y_out_double_2_7_axb_10),.CI(Y_out_double_2_7_cry_9),.O(Y_out_double_2_7[10:10]));
  MUXCY_L Y_out_double_2_7_cry_10_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_9),.S(Y_out_double_2_7_axb_10),.LO(Y_out_double_2_7_cry_10));
  XORCY Y_out_double_2_7_s_9(.LI(Y_out_double_2_7_axb_9),.CI(Y_out_double_2_7_cry_8),.O(Y_out_double_2_7[9:9]));
  MUXCY_L Y_out_double_2_7_cry_9_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_8),.S(Y_out_double_2_7_axb_9),.LO(Y_out_double_2_7_cry_9));
  XORCY Y_out_double_2_7_s_8(.LI(Y_out_double_2_7_axb_8),.CI(Y_out_double_2_7_cry_7),.O(Y_out_double_2_7[8:8]));
  MUXCY_L Y_out_double_2_7_cry_8_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_7),.S(Y_out_double_2_7_axb_8),.LO(Y_out_double_2_7_cry_8));
  XORCY Y_out_double_2_7_s_7(.LI(Y_out_double_2_7_axb_7),.CI(Y_out_double_2_7_cry_6),.O(Y_out_double_2_7[7:7]));
  MUXCY_L Y_out_double_2_7_cry_7_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_6),.S(Y_out_double_2_7_axb_7),.LO(Y_out_double_2_7_cry_7));
  XORCY Y_out_double_2_7_s_6(.LI(Y_out_double_2_7_axb_6),.CI(Y_out_double_2_7_cry_5),.O(Y_out_double_2_7[6:6]));
  MUXCY_L Y_out_double_2_7_cry_6_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_5),.S(Y_out_double_2_7_axb_6),.LO(Y_out_double_2_7_cry_6));
  XORCY Y_out_double_2_7_s_5(.LI(Y_out_double_2_7_axb_5),.CI(Y_out_double_2_7_cry_4),.O(Y_out_double_2_7[5:5]));
  MUXCY_L Y_out_double_2_7_cry_5_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_4),.S(Y_out_double_2_7_axb_5),.LO(Y_out_double_2_7_cry_5));
  XORCY Y_out_double_2_7_s_4(.LI(Y_out_double_2_7_axb_4),.CI(Y_out_double_2_7_cry_3),.O(Y_out_double_2_7[4:4]));
  MUXCY_L Y_out_double_2_7_cry_4_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_3),.S(Y_out_double_2_7_axb_4),.LO(Y_out_double_2_7_cry_4));
  XORCY Y_out_double_2_7_s_3(.LI(Y_out_double_2_7_axb_3),.CI(Y_out_double_2_7_cry_2),.O(Y_out_double_2_7[3:3]));
  MUXCY_L Y_out_double_2_7_cry_3_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_2),.S(Y_out_double_2_7_axb_3),.LO(Y_out_double_2_7_cry_3));
  XORCY Y_out_double_2_7_s_2(.LI(Y_out_double_2_7_axb_2),.CI(Y_out_double_2_7_cry_1),.O(Y_out_double_2_7[2:2]));
  MUXCY_L Y_out_double_2_7_cry_2_cZ(.DI(GND),.CI(Y_out_double_2_7_cry_1),.S(Y_out_double_2_7_axb_2),.LO(Y_out_double_2_7_cry_2));
  MUXCY_L Y_out_double_2_7_cry_1_cZ(.DI(VCC),.CI(GND),.S(pgZFF_X0_i[1:1]),.LO(Y_out_double_2_7_cry_1));
  XORCY Y_out_double_2_s_17(.LI(Y_out_double_2_axb_17),.CI(Y_out_double_2_cry_16),.O(Y_out_double_2[17:17]));
  XORCY Y_out_double_2_s_16(.LI(Y_out_double_2_axb_16),.CI(Y_out_double_2_cry_15),.O(Y_out_double_2[16:16]));
  MUXCY_L Y_out_double_2_cry_16_cZ(.DI(Y_out_double_2_4[16:16]),.CI(Y_out_double_2_cry_15),.S(Y_out_double_2_axb_16),.LO(Y_out_double_2_cry_16));
  XORCY Y_out_double_2_s_15(.LI(Y_out_double_2_axb_15),.CI(Y_out_double_2_cry_14),.O(Y_out_double_2[15:15]));
  MUXCY_L Y_out_double_2_cry_15_cZ(.DI(Y_out_double_2_4[15:15]),.CI(Y_out_double_2_cry_14),.S(Y_out_double_2_axb_15),.LO(Y_out_double_2_cry_15));
  XORCY Y_out_double_2_s_14(.LI(Y_out_double_2_axb_14),.CI(Y_out_double_2_cry_13),.O(Y_out_double_2[14:14]));
  MUXCY_L Y_out_double_2_cry_14_cZ(.DI(Y_out_double_2_4[14:14]),.CI(Y_out_double_2_cry_13),.S(Y_out_double_2_axb_14),.LO(Y_out_double_2_cry_14));
  XORCY Y_out_double_2_s_13(.LI(Y_out_double_2_axb_13),.CI(Y_out_double_2_cry_12),.O(Y_out_double_2[13:13]));
  MUXCY_L Y_out_double_2_cry_13_cZ(.DI(Y_out_double_2_4[13:13]),.CI(Y_out_double_2_cry_12),.S(Y_out_double_2_axb_13),.LO(Y_out_double_2_cry_13));
  XORCY Y_out_double_2_s_12(.LI(Y_out_double_2_axb_12),.CI(Y_out_double_2_cry_11),.O(Y_out_double_2[12:12]));
  MUXCY_L Y_out_double_2_cry_12_cZ(.DI(Y_out_double_2_4[12:12]),.CI(Y_out_double_2_cry_11),.S(Y_out_double_2_axb_12),.LO(Y_out_double_2_cry_12));
  XORCY Y_out_double_2_s_11(.LI(Y_out_double_2_axb_11),.CI(Y_out_double_2_cry_10),.O(Y_out_double_2[11:11]));
  MUXCY_L Y_out_double_2_cry_11_cZ(.DI(Y_out_double_2_4[11:11]),.CI(Y_out_double_2_cry_10),.S(Y_out_double_2_axb_11),.LO(Y_out_double_2_cry_11));
  XORCY Y_out_double_2_s_10(.LI(Y_out_double_2_axb_10),.CI(Y_out_double_2_cry_9),.O(Y_out_double_2[10:10]));
  MUXCY_L Y_out_double_2_cry_10_cZ(.DI(Y_out_double_2_4[10:10]),.CI(Y_out_double_2_cry_9),.S(Y_out_double_2_axb_10),.LO(Y_out_double_2_cry_10));
  XORCY Y_out_double_2_s_9(.LI(Y_out_double_2_axb_9),.CI(Y_out_double_2_cry_8),.O(Y_out_double_2[9:9]));
  MUXCY_L Y_out_double_2_cry_9_cZ(.DI(Y_out_double_2_4[9:9]),.CI(Y_out_double_2_cry_8),.S(Y_out_double_2_axb_9),.LO(Y_out_double_2_cry_9));
  XORCY Y_out_double_2_s_8(.LI(Y_out_double_2_axb_8),.CI(Y_out_double_2_cry_7),.O(Y_out_double_2[8:8]));
  MUXCY_L Y_out_double_2_cry_8_cZ(.DI(Y_out_double_2_4[8:8]),.CI(Y_out_double_2_cry_7),.S(Y_out_double_2_axb_8),.LO(Y_out_double_2_cry_8));
  XORCY Y_out_double_2_s_7(.LI(Y_out_double_2_axb_7),.CI(Y_out_double_2_cry_6),.O(Y_out_double_2[7:7]));
  MUXCY_L Y_out_double_2_cry_7_cZ(.DI(Y_out_double_2_4[7:7]),.CI(Y_out_double_2_cry_6),.S(Y_out_double_2_axb_7),.LO(Y_out_double_2_cry_7));
  XORCY Y_out_double_2_s_6(.LI(Y_out_double_2_axb_6),.CI(Y_out_double_2_cry_5),.O(Y_out_double_2[6:6]));
  MUXCY_L Y_out_double_2_cry_6_cZ(.DI(Y_out_double_2_4[6:6]),.CI(Y_out_double_2_cry_5),.S(Y_out_double_2_axb_6),.LO(Y_out_double_2_cry_6));
  XORCY Y_out_double_2_s_5(.LI(Y_out_double_2_axb_5),.CI(Y_out_double_2_cry_4),.O(Y_out_double_2[5:5]));
  MUXCY_L Y_out_double_2_cry_5_cZ(.DI(Y_out_double_2_4[5:5]),.CI(Y_out_double_2_cry_4),.S(Y_out_double_2_axb_5),.LO(Y_out_double_2_cry_5));
  XORCY Y_out_double_2_s_4(.LI(Y_out_double_2_axb_4),.CI(Y_out_double_2_cry_3),.O(Y_out_double_2[4:4]));
  MUXCY_L Y_out_double_2_cry_4_cZ(.DI(Y_out_double_2_4[4:4]),.CI(Y_out_double_2_cry_3),.S(Y_out_double_2_axb_4),.LO(Y_out_double_2_cry_4));
  XORCY Y_out_double_2_s_3(.LI(Y_out_double_2_axb_3),.CI(Y_out_double_2_cry_2),.O(Y_out_double_2[3:3]));
  MUXCY_L Y_out_double_2_cry_3_cZ(.DI(Y_out_double_2_4[3:3]),.CI(Y_out_double_2_cry_2),.S(Y_out_double_2_axb_3),.LO(Y_out_double_2_cry_3));
  XORCY Y_out_double_2_s_2(.LI(Y_out_double_2_axb_2),.CI(Y_out_double_2_cry_1),.O(Y_out_double_2[2:2]));
  MUXCY_L Y_out_double_2_cry_2_cZ(.DI(Y_out_double_2_4[2:2]),.CI(Y_out_double_2_cry_1),.S(Y_out_double_2_axb_2),.LO(Y_out_double_2_cry_2));
  XORCY Y_out_double_2_s_1(.LI(Y_out_double_2_axb_1),.CI(Y_out_double_2_cry_0),.O(Y_out_double_2[1:1]));
  MUXCY_L Y_out_double_2_cry_1_cZ(.DI(Y_out_double_2_4[1:1]),.CI(Y_out_double_2_cry_0),.S(Y_out_double_2_axb_1),.LO(Y_out_double_2_cry_1));
  MUXCY_L Y_out_double_2_cry_0_cZ(.DI(Y_out_double_2_4[0:0]),.CI(GND),.S(Y_out_double_2[0:0]),.LO(Y_out_double_2_cry_0));
  XORCY un10_8_s_28(.LI(un10_8_axb_28),.CI(un10_8_cry_27),.O(un10_8[47:47]));
  XORCY un10_8_s_27(.LI(un10_8_axb_27),.CI(un10_8_cry_26),.O(un10_8[45:45]));
  MUXCY_L un10_8_cry_27_cZ(.DI(GND),.CI(un10_8_cry_26),.S(un10_8_axb_27),.LO(un10_8_cry_27));
  XORCY un10_8_s_26(.LI(un10_8_axb_26),.CI(un10_8_cry_25),.O(un10_8[44:44]));
  MUXCY_L un10_8_cry_26_cZ(.DI(GND),.CI(un10_8_cry_25),.S(un10_8_axb_26),.LO(un10_8_cry_26));
  XORCY un10_8_s_25(.LI(un10_8_axb_25),.CI(un10_8_cry_24),.O(un10_8[43:43]));
  MUXCY_L un10_8_cry_25_cZ(.DI(ZFF_Y2[15:15]),.CI(un10_8_cry_24),.S(un10_8_axb_25),.LO(un10_8_cry_25));
  XORCY un10_8_s_24(.LI(un10_8_axb_24),.CI(un10_8_cry_23),.O(un10_8[42:42]));
  MUXCY_L un10_8_cry_24_cZ(.DI(un10_8_o5_23),.CI(un10_8_cry_23),.S(un10_8_axb_24),.LO(un10_8_cry_24));
  XORCY un10_8_s_23(.LI(un10_8_axb_23),.CI(un10_8_cry_22),.O(un10_8[41:41]));
  MUXCY_L un10_8_cry_23_cZ(.DI(un10_8_o5_22),.CI(un10_8_cry_22),.S(un10_8_axb_23),.LO(un10_8_cry_23));
  XORCY un10_8_s_22(.LI(un10_8_axb_22),.CI(un10_8_cry_21),.O(un10_8[40:40]));
  MUXCY_L un10_8_cry_22_cZ(.DI(un10_8_o5_21),.CI(un10_8_cry_21),.S(un10_8_axb_22),.LO(un10_8_cry_22));
  XORCY un10_8_s_21(.LI(un10_8_axb_21),.CI(un10_8_cry_20),.O(un10_8[39:39]));
  MUXCY_L un10_8_cry_21_cZ(.DI(un10_8_o5_20),.CI(un10_8_cry_20),.S(un10_8_axb_21),.LO(un10_8_cry_21));
  XORCY un10_8_s_20(.LI(un10_8_axb_20),.CI(un10_8_cry_19),.O(un10_8[38:38]));
  MUXCY_L un10_8_cry_20_cZ(.DI(un10_8_o5_19),.CI(un10_8_cry_19),.S(un10_8_axb_20),.LO(un10_8_cry_20));
  XORCY un10_8_s_19(.LI(un10_8_axb_19),.CI(un10_8_cry_18),.O(un10_8[37:37]));
  MUXCY_L un10_8_cry_19_cZ(.DI(un10_8_o5_18),.CI(un10_8_cry_18),.S(un10_8_axb_19),.LO(un10_8_cry_19));
  XORCY un10_8_s_18(.LI(un10_8_axb_18),.CI(un10_8_cry_17),.O(un10_8[36:36]));
  MUXCY_L un10_8_cry_18_cZ(.DI(un10_8_o5_17),.CI(un10_8_cry_17),.S(un10_8_axb_18),.LO(un10_8_cry_18));
  XORCY un10_8_s_17(.LI(un10_8_axb_17),.CI(un10_8_cry_16),.O(un10_8[35:35]));
  MUXCY_L un10_8_cry_17_cZ(.DI(un10_8_o5_16),.CI(un10_8_cry_16),.S(un10_8_axb_17),.LO(un10_8_cry_17));
  XORCY un10_8_s_16(.LI(un10_8_axb_16),.CI(un10_8_cry_15),.O(un10_8[34:34]));
  MUXCY_L un10_8_cry_16_cZ(.DI(un10_8_o5_15),.CI(un10_8_cry_15),.S(un10_8_axb_16),.LO(un10_8_cry_16));
  XORCY un10_8_s_15(.LI(un10_8_axb_15),.CI(un10_8_cry_14),.O(un10_8[33:33]));
  MUXCY_L un10_8_cry_15_cZ(.DI(un10_8_o5_14),.CI(un10_8_cry_14),.S(un10_8_axb_15),.LO(un10_8_cry_15));
  XORCY un10_8_s_14(.LI(un10_8_axb_14),.CI(un10_8_cry_13),.O(un10_8[32:32]));
  MUXCY_L un10_8_cry_14_cZ(.DI(un10_8_o5_13),.CI(un10_8_cry_13),.S(un10_8_axb_14),.LO(un10_8_cry_14));
  XORCY un10_8_s_13(.LI(un10_8_axb_13),.CI(un10_8_cry_12),.O(un10_8[31:31]));
  MUXCY_L un10_8_cry_13_cZ(.DI(un10_8_o5_12),.CI(un10_8_cry_12),.S(un10_8_axb_13),.LO(un10_8_cry_13));
  XORCY un10_8_s_12(.LI(un10_8_axb_12),.CI(un10_8_cry_11),.O(un10_8[30:30]));
  MUXCY_L un10_8_cry_12_cZ(.DI(un10_8_o5_11),.CI(un10_8_cry_11),.S(un10_8_axb_12),.LO(un10_8_cry_12));
  XORCY un10_8_s_11(.LI(un10_8_axb_11),.CI(un10_8_cry_10),.O(un10_8[29:29]));
  MUXCY_L un10_8_cry_11_cZ(.DI(un10_8_cry_11_RNO),.CI(un10_8_cry_10),.S(un10_8_axb_11),.LO(un10_8_cry_11));
  XORCY un10_8_s_10(.LI(un10_8_axb_10),.CI(un10_8_cry_9),.O(un10_8[28:28]));
  MUXCY_L un10_8_cry_10_cZ(.DI(N_2973_i),.CI(un10_8_cry_9),.S(un10_8_axb_10),.LO(un10_8_cry_10));
  XORCY un10_8_s_9(.LI(un10_8_axb_9),.CI(un10_8_cry_8),.O(un10_8[27:27]));
  MUXCY_L un10_8_cry_9_cZ(.DI(ZFF_Y2[1:1]),.CI(un10_8_cry_8),.S(un10_8_axb_9),.LO(un10_8_cry_9));
  XORCY un10_8_s_8(.LI(un10_8_axb_8),.CI(un10_8_cry_7),.O(un10_8[26:26]));
  MUXCY_L un10_8_cry_8_cZ(.DI(ZFF_Y2[0:0]),.CI(un10_8_cry_7),.S(un10_8_axb_8),.LO(un10_8_cry_8));
  XORCY un10_8_s_7(.LI(un10_8_axb_7),.CI(un10_8_cry_6),.O(un10_8[25:25]));
  MUXCY_L un10_8_cry_7_cZ(.DI(GND),.CI(un10_8_cry_6),.S(un10_8_axb_7),.LO(un10_8_cry_7));
  XORCY un10_8_s_6(.LI(un10_8_axb_6),.CI(un10_8_cry_5),.O(un10_8[24:24]));
  MUXCY_L un10_8_cry_6_cZ(.DI(GND),.CI(un10_8_cry_5),.S(un10_8_axb_6),.LO(un10_8_cry_6));
  XORCY un10_8_s_5(.LI(un10_8_axb_5),.CI(un10_8_cry_4),.O(un10_8[23:23]));
  MUXCY_L un10_8_cry_5_cZ(.DI(GND),.CI(un10_8_cry_4),.S(un10_8_axb_5),.LO(un10_8_cry_5));
  XORCY un10_8_s_4(.LI(un10_8_axb_4),.CI(un10_8_cry_3),.O(un10_8[22:22]));
  MUXCY_L un10_8_cry_4_cZ(.DI(ZFF_Y2_fast[17:17]),.CI(un10_8_cry_3),.S(un10_8_axb_4),.LO(un10_8_cry_4));
  XORCY un10_8_s_3(.LI(un10_8_axb_3),.CI(un10_8_cry_2),.O(un10_8[21:21]));
  MUXCY_L un10_8_cry_3_cZ(.DI(ZFF_Y2_fast[17:17]),.CI(un10_8_cry_2),.S(un10_8_axb_3),.LO(un10_8_cry_3));
  XORCY un10_8_s_2(.LI(un10_8_axb_2),.CI(un10_8_cry_1),.O(un10_8[20:20]));
  MUXCY_L un10_8_cry_2_cZ(.DI(ZFF_Y2_fast[17:17]),.CI(un10_8_cry_1),.S(un10_8_axb_2),.LO(un10_8_cry_2));
  XORCY un10_8_s_1(.LI(un10_8_axb_1),.CI(un10_8_cry_0),.O(un10_8[19:19]));
  MUXCY_L un10_8_cry_1_cZ(.DI(ZFF_Y2_fast[17:17]),.CI(un10_8_cry_0),.S(un10_8_axb_1),.LO(un10_8_cry_1));
  XORCY un10_8_s_0(.LI(un10_8_axb_0),.CI(un10_8_cry_0_cy),.O(un10_8[18:18]));
  MUXCY_L un10_8_cry_0_cZ(.DI(ZFF_Y2_fast[17:17]),.CI(un10_8_cry_0_cy),.S(un10_8_axb_0),.LO(un10_8_cry_0));
  XORCY un8_0_8_s_26(.LI(un8_0_8_axb_26),.CI(un8_0_8_cry_25),.O(un8_0_8[36:36]));
  MUXCY_L un8_0_8_cry_26(.DI(ZFF_X2[15:15]),.CI(un8_0_8_cry_25),.S(un8_0_8_axb_26),.LO(un8_0_8[38:38]));
  XORCY un8_0_8_s_25(.LI(un8_0_8_axb_25),.CI(un8_0_8_cry_24),.O(un8_0_8[35:35]));
  MUXCY_L un8_0_8_cry_25_cZ(.DI(ZFF_X2[14:14]),.CI(un8_0_8_cry_24),.S(un8_0_8_axb_25),.LO(un8_0_8_cry_25));
  XORCY un8_0_8_s_24(.LI(un8_0_8_axb_24),.CI(un8_0_8_cry_23),.O(un8_0_8[34:34]));
  MUXCY_L un8_0_8_cry_24_cZ(.DI(ZFF_X2[13:13]),.CI(un8_0_8_cry_23),.S(un8_0_8_axb_24),.LO(un8_0_8_cry_24));
  XORCY un8_0_8_s_23(.LI(un8_0_8_axb_23),.CI(un8_0_8_cry_22),.O(un8_0_8[33:33]));
  MUXCY_L un8_0_8_cry_23_cZ(.DI(ZFF_X2[12:12]),.CI(un8_0_8_cry_22),.S(un8_0_8_axb_23),.LO(un8_0_8_cry_23));
  XORCY un8_0_8_s_22(.LI(un8_0_8_axb_22),.CI(un8_0_8_cry_21),.O(un8_0_8[32:32]));
  MUXCY_L un8_0_8_cry_22_cZ(.DI(ZFF_X2[11:11]),.CI(un8_0_8_cry_21),.S(un8_0_8_axb_22),.LO(un8_0_8_cry_22));
  XORCY un8_0_8_s_21(.LI(un8_0_8_axb_21),.CI(un8_0_8_cry_20),.O(un8_0_8[31:31]));
  MUXCY_L un8_0_8_cry_21_cZ(.DI(N_3180_i),.CI(un8_0_8_cry_20),.S(un8_0_8_axb_21),.LO(un8_0_8_cry_21));
  XORCY un8_0_8_s_20(.LI(un8_0_8_axb_20),.CI(un8_0_8_cry_19),.O(un8_0_8[30:30]));
  MUXCY_L un8_0_8_cry_20_cZ(.DI(un8_0_8_cry_20_RNO),.CI(un8_0_8_cry_19),.S(un8_0_8_axb_20),.LO(un8_0_8_cry_20));
  XORCY un8_0_8_s_19(.LI(un8_0_8_axb_19),.CI(un8_0_8_cry_18),.O(un8_0_8[29:29]));
  MUXCY_L un8_0_8_cry_19_cZ(.DI(un8_0_8_cry_19_RNO),.CI(un8_0_8_cry_18),.S(un8_0_8_axb_19),.LO(un8_0_8_cry_19));
  XORCY un8_0_8_s_18(.LI(un8_0_8_axb_18),.CI(un8_0_8_cry_17),.O(un8_0_8[28:28]));
  MUXCY_L un8_0_8_cry_18_cZ(.DI(un8_0_8_cry_18_RNO),.CI(un8_0_8_cry_17),.S(un8_0_8_axb_18),.LO(un8_0_8_cry_18));
  XORCY un8_0_8_s_17(.LI(un8_0_8_axb_17),.CI(un8_0_8_cry_16),.O(un8_0_8[27:27]));
  MUXCY_L un8_0_8_cry_17_cZ(.DI(un8_0_8_cry_17_RNO),.CI(un8_0_8_cry_16),.S(un8_0_8_axb_17),.LO(un8_0_8_cry_17));
  XORCY un8_0_8_s_16(.LI(un8_0_8_axb_16),.CI(un8_0_8_cry_15),.O(un8_0_8[26:26]));
  MUXCY_L un8_0_8_cry_16_cZ(.DI(un8_0_8_cry_16_RNO),.CI(un8_0_8_cry_15),.S(un8_0_8_axb_16),.LO(un8_0_8_cry_16));
  XORCY un8_0_8_s_15(.LI(un8_0_8_axb_15),.CI(un8_0_8_cry_14),.O(un8_0_8[25:25]));
  MUXCY_L un8_0_8_cry_15_cZ(.DI(un8_0_6_1_scalar),.CI(un8_0_8_cry_14),.S(un8_0_8_axb_15),.LO(un8_0_8_cry_15));
  XORCY un8_0_8_s_14(.LI(un8_0_8_axb_14),.CI(un8_0_8_cry_13),.O(un8_0_8[24:24]));
  MUXCY_L un8_0_8_cry_14_cZ(.DI(un8_0_8_cry_14_RNO),.CI(un8_0_8_cry_13),.S(un8_0_8_axb_14),.LO(un8_0_8_cry_14));
  XORCY un8_0_8_s_13(.LI(un8_0_8_axb_13),.CI(un8_0_8_cry_12),.O(un8_0_8[23:23]));
  MUXCY_L un8_0_8_cry_13_cZ(.DI(un8_0_8_cry_13_RNO),.CI(un8_0_8_cry_12),.S(un8_0_8_axb_13),.LO(un8_0_8_cry_13));
  XORCY un8_0_8_s_12(.LI(un8_0_8_axb_12),.CI(un8_0_8_cry_11),.O(un8_0_8[22:22]));
  MUXCY_L un8_0_8_cry_12_cZ(.DI(un8_0_8_o5_11),.CI(un8_0_8_cry_11),.S(un8_0_8_axb_12),.LO(un8_0_8_cry_12));
  XORCY un8_0_8_s_11(.LI(un8_0_8_axb_11),.CI(un8_0_8_cry_10),.O(un8_0_8[21:21]));
  MUXCY_L un8_0_8_cry_11_cZ(.DI(un8_0_8_o5_10),.CI(un8_0_8_cry_10),.S(un8_0_8_axb_11),.LO(un8_0_8_cry_11));
  XORCY un8_0_8_s_10(.LI(un8_0_8_axb_10),.CI(un8_0_8_cry_9),.O(un8_0_8[20:20]));
  MUXCY_L un8_0_8_cry_10_cZ(.DI(un8_0_8_cry_10_RNO),.CI(un8_0_8_cry_9),.S(un8_0_8_axb_10),.LO(un8_0_8_cry_10));
  XORCY un8_0_8_s_9(.LI(un8_0_8_axb_9),.CI(un8_0_8_cry_8),.O(un8_0_8[19:19]));
  MUXCY_L un8_0_8_cry_9_cZ(.DI(un8_0_8_cry_9_RNO),.CI(un8_0_8_cry_8),.S(un8_0_8_axb_9),.LO(un8_0_8_cry_9));
  XORCY un8_0_8_s_8(.LI(un8_0_8_axb_8),.CI(un8_0_8_cry_7),.O(un8_0_8[18:18]));
  MUXCY_L un8_0_8_cry_8_cZ(.DI(un8_0_8_cry_8_RNO),.CI(un8_0_8_cry_7),.S(un8_0_8_axb_8),.LO(un8_0_8_cry_8));
  XORCY un8_0_8_s_7(.LI(un8_0_8_axb_7),.CI(un8_0_8_cry_6),.O(un8_0_8[17:17]));
  MUXCY_L un8_0_8_cry_7_cZ(.DI(un8_0_8_cry_7_RNO),.CI(un8_0_8_cry_6),.S(un8_0_8_axb_7),.LO(un8_0_8_cry_7));
  XORCY un8_0_8_s_6(.LI(un8_0_8_axb_6),.CI(un8_0_8_cry_5),.O(un8_0_8[16:16]));
  MUXCY_L un8_0_8_cry_6_cZ(.DI(un8_0_8_cry_6_RNO),.CI(un8_0_8_cry_5),.S(un8_0_8_axb_6),.LO(un8_0_8_cry_6));
  XORCY un8_0_8_s_5(.LI(un8_0_8_axb_5),.CI(un8_0_8_cry_4),.O(un8_0_8[15:15]));
  MUXCY_L un8_0_8_cry_5_cZ(.DI(un8_0_8_o5_4),.CI(un8_0_8_cry_4),.S(un8_0_8_axb_5),.LO(un8_0_8_cry_5));
  XORCY un8_0_8_s_4(.LI(un8_0_8_axb_4),.CI(un8_0_8_cry_3),.O(un8_0_8[14:14]));
  MUXCY_L un8_0_8_cry_4_cZ(.DI(un8_0_8_cry_4_RNO),.CI(un8_0_8_cry_3),.S(un8_0_8_axb_4),.LO(un8_0_8_cry_4));
  XORCY un8_0_8_s_3(.LI(un8_0_8_axb_3),.CI(un8_0_8_cry_2),.O(un8_0_8[13:13]));
  MUXCY_L un8_0_8_cry_3_cZ(.DI(un8_0_8_cry_3_RNO),.CI(un8_0_8_cry_2),.S(un8_0_8_axb_3),.LO(un8_0_8_cry_3));
  XORCY un8_0_8_s_2(.LI(un8_0_8_axb_2),.CI(un8_0_8_cry_1),.O(un8_0_8[12:12]));
  MUXCY_L un8_0_8_cry_2_cZ(.DI(GND),.CI(un8_0_8_cry_1),.S(un8_0_8_axb_2),.LO(un8_0_8_cry_2));
  XORCY un8_0_8_s_1(.LI(un8_0_8_axb_1),.CI(un8_0_8_cry_0),.O(un8_0_8[11:11]));
  MUXCY_L un8_0_8_cry_1_cZ(.DI(ZFF_X2_3_rep1),.CI(un8_0_8_cry_0),.S(un8_0_8_axb_1),.LO(un8_0_8_cry_1));
  MUXCY_L un8_0_8_cry_0_cZ(.DI(ZFF_X2_fast[2:2]),.CI(GND),.S(un8_0_8[10:10]),.LO(un8_0_8_cry_0));
  XORCY un6_0_8_s_26(.LI(un6_0_8_axb_26),.CI(un6_0_8_cry_25),.O(un6_0_8[36:36]));
  MUXCY_L un6_0_8_cry_26(.DI(ZFF_X0[15:15]),.CI(un6_0_8_cry_25),.S(un6_0_8_axb_26),.LO(un6_0_8[38:38]));
  XORCY un6_0_8_s_25(.LI(un6_0_8_axb_25),.CI(un6_0_8_cry_24),.O(un6_0_8[35:35]));
  MUXCY_L un6_0_8_cry_25_cZ(.DI(ZFF_X0[14:14]),.CI(un6_0_8_cry_24),.S(un6_0_8_axb_25),.LO(un6_0_8_cry_25));
  XORCY un6_0_8_s_24(.LI(un6_0_8_axb_24),.CI(un6_0_8_cry_23),.O(un6_0_8[34:34]));
  MUXCY_L un6_0_8_cry_24_cZ(.DI(ZFF_X0[13:13]),.CI(un6_0_8_cry_23),.S(un6_0_8_axb_24),.LO(un6_0_8_cry_24));
  XORCY un6_0_8_s_23(.LI(un6_0_8_axb_23),.CI(un6_0_8_cry_22),.O(un6_0_8[33:33]));
  MUXCY_L un6_0_8_cry_23_cZ(.DI(ZFF_X0[12:12]),.CI(un6_0_8_cry_22),.S(un6_0_8_axb_23),.LO(un6_0_8_cry_23));
  XORCY un6_0_8_s_22(.LI(un6_0_8_axb_22),.CI(un6_0_8_cry_21),.O(un6_0_8[32:32]));
  MUXCY_L un6_0_8_cry_22_cZ(.DI(ZFF_X0[11:11]),.CI(un6_0_8_cry_21),.S(un6_0_8_axb_22),.LO(un6_0_8_cry_22));
  XORCY un6_0_8_s_21(.LI(un6_0_8_axb_21),.CI(un6_0_8_cry_20),.O(un6_0_8[31:31]));
  MUXCY_L un6_0_8_cry_21_cZ(.DI(N_2366_i),.CI(un6_0_8_cry_20),.S(un6_0_8_axb_21),.LO(un6_0_8_cry_21));
  XORCY un6_0_8_s_20(.LI(un6_0_8_axb_20),.CI(un6_0_8_cry_19),.O(un6_0_8[30:30]));
  MUXCY_L un6_0_8_cry_20_cZ(.DI(un6_0_8_cry_20_RNO),.CI(un6_0_8_cry_19),.S(un6_0_8_axb_20),.LO(un6_0_8_cry_20));
  XORCY un6_0_8_s_19(.LI(un6_0_8_axb_19),.CI(un6_0_8_cry_18),.O(un6_0_8[29:29]));
  MUXCY_L un6_0_8_cry_19_cZ(.DI(un6_0_8_cry_19_RNO),.CI(un6_0_8_cry_18),.S(un6_0_8_axb_19),.LO(un6_0_8_cry_19));
  XORCY un6_0_8_s_18(.LI(un6_0_8_axb_18),.CI(un6_0_8_cry_17),.O(un6_0_8[28:28]));
  MUXCY_L un6_0_8_cry_18_cZ(.DI(un6_0_8_cry_18_RNO),.CI(un6_0_8_cry_17),.S(un6_0_8_axb_18),.LO(un6_0_8_cry_18));
  XORCY un6_0_8_s_17(.LI(un6_0_8_axb_17),.CI(un6_0_8_cry_16),.O(un6_0_8[27:27]));
  MUXCY_L un6_0_8_cry_17_cZ(.DI(un6_0_8_cry_17_RNO),.CI(un6_0_8_cry_16),.S(un6_0_8_axb_17),.LO(un6_0_8_cry_17));
  XORCY un6_0_8_s_16(.LI(un6_0_8_axb_16),.CI(un6_0_8_cry_15),.O(un6_0_8[26:26]));
  MUXCY_L un6_0_8_cry_16_cZ(.DI(un6_0_8_cry_16_RNO),.CI(un6_0_8_cry_15),.S(un6_0_8_axb_16),.LO(un6_0_8_cry_16));
  XORCY un6_0_8_s_15(.LI(un6_0_8_axb_15),.CI(un6_0_8_cry_14),.O(un6_0_8[25:25]));
  MUXCY_L un6_0_8_cry_15_cZ(.DI(un6_0_6_1_scalar),.CI(un6_0_8_cry_14),.S(un6_0_8_axb_15),.LO(un6_0_8_cry_15));
  XORCY un6_0_8_s_14(.LI(un6_0_8_axb_14),.CI(un6_0_8_cry_13),.O(un6_0_8[24:24]));
  MUXCY_L un6_0_8_cry_14_cZ(.DI(un6_0_8_cry_14_RNO),.CI(un6_0_8_cry_13),.S(un6_0_8_axb_14),.LO(un6_0_8_cry_14));
  XORCY un6_0_8_s_13(.LI(un6_0_8_axb_13),.CI(un6_0_8_cry_12),.O(un6_0_8[23:23]));
  MUXCY_L un6_0_8_cry_13_cZ(.DI(un6_0_8_cry_13_RNO),.CI(un6_0_8_cry_12),.S(un6_0_8_axb_13),.LO(un6_0_8_cry_13));
  XORCY un6_0_8_s_12(.LI(un6_0_8_axb_12),.CI(un6_0_8_cry_11),.O(un6_0_8[22:22]));
  MUXCY_L un6_0_8_cry_12_cZ(.DI(un6_0_8_o5_11),.CI(un6_0_8_cry_11),.S(un6_0_8_axb_12),.LO(un6_0_8_cry_12));
  XORCY un6_0_8_s_11(.LI(un6_0_8_axb_11),.CI(un6_0_8_cry_10),.O(un6_0_8[21:21]));
  MUXCY_L un6_0_8_cry_11_cZ(.DI(un6_0_8_o5_10),.CI(un6_0_8_cry_10),.S(un6_0_8_axb_11),.LO(un6_0_8_cry_11));
  XORCY un6_0_8_s_10(.LI(un6_0_8_axb_10),.CI(un6_0_8_cry_9),.O(un6_0_8[20:20]));
  MUXCY_L un6_0_8_cry_10_cZ(.DI(un6_0_8_cry_10_RNO),.CI(un6_0_8_cry_9),.S(un6_0_8_axb_10),.LO(un6_0_8_cry_10));
  XORCY un6_0_8_s_9(.LI(un6_0_8_axb_9),.CI(un6_0_8_cry_8),.O(un6_0_8[19:19]));
  MUXCY_L un6_0_8_cry_9_cZ(.DI(un6_0_8_cry_9_RNO),.CI(un6_0_8_cry_8),.S(un6_0_8_axb_9),.LO(un6_0_8_cry_9));
  XORCY un6_0_8_s_8(.LI(un6_0_8_axb_8),.CI(un6_0_8_cry_7),.O(un6_0_8[18:18]));
  MUXCY_L un6_0_8_cry_8_cZ(.DI(un6_0_8_cry_8_RNO),.CI(un6_0_8_cry_7),.S(un6_0_8_axb_8),.LO(un6_0_8_cry_8));
  XORCY un6_0_8_s_7(.LI(un6_0_8_axb_7),.CI(un6_0_8_cry_6),.O(un6_0_8[17:17]));
  MUXCY_L un6_0_8_cry_7_cZ(.DI(un6_0_8_cry_7_RNO),.CI(un6_0_8_cry_6),.S(un6_0_8_axb_7),.LO(un6_0_8_cry_7));
  XORCY un6_0_8_s_6(.LI(un6_0_8_axb_6),.CI(un6_0_8_cry_5),.O(un6_0_8[16:16]));
  MUXCY_L un6_0_8_cry_6_cZ(.DI(un6_0_8_cry_6_RNO),.CI(un6_0_8_cry_5),.S(un6_0_8_axb_6),.LO(un6_0_8_cry_6));
  XORCY un6_0_8_s_5(.LI(un6_0_8_axb_5),.CI(un6_0_8_cry_4),.O(un6_0_8[15:15]));
  MUXCY_L un6_0_8_cry_5_cZ(.DI(un6_0_8_o5_4),.CI(un6_0_8_cry_4),.S(un6_0_8_axb_5),.LO(un6_0_8_cry_5));
  XORCY un6_0_8_s_4(.LI(un6_0_8_axb_4),.CI(un6_0_8_cry_3),.O(un6_0_8[14:14]));
  MUXCY_L un6_0_8_cry_4_cZ(.DI(un6_0_8_cry_4_RNO),.CI(un6_0_8_cry_3),.S(un6_0_8_axb_4),.LO(un6_0_8_cry_4));
  XORCY un6_0_8_s_3(.LI(un6_0_8_axb_3),.CI(un6_0_8_cry_2),.O(un6_0_8[13:13]));
  MUXCY_L un6_0_8_cry_3_cZ(.DI(un6_0_8_cry_3_RNO),.CI(un6_0_8_cry_2),.S(un6_0_8_axb_3),.LO(un6_0_8_cry_3));
  XORCY un6_0_8_s_2(.LI(un6_0_8_axb_2),.CI(un6_0_8_cry_1),.O(un6_0_8[12:12]));
  MUXCY_L un6_0_8_cry_2_cZ(.DI(GND),.CI(un6_0_8_cry_1),.S(un6_0_8_axb_2),.LO(un6_0_8_cry_2));
  XORCY un6_0_8_s_1(.LI(un6_0_8_axb_1),.CI(un6_0_8_cry_0),.O(un6_0_8[11:11]));
  MUXCY_L un6_0_8_cry_1_cZ(.DI(ZFF_X0_3_rep1),.CI(un6_0_8_cry_0),.S(un6_0_8_axb_1),.LO(un6_0_8_cry_1));
  MUXCY_L un6_0_8_cry_0_cZ(.DI(ZFF_X0_fast[2:2]),.CI(GND),.S(un6_0_8[10:10]),.LO(un6_0_8_cry_0));
  XORCY un7_0_8_s_28(.LI(un7_0_8_axb_28),.CI(un7_0_8_cry_27),.O(un7_0_8[37:37]));
  MUXCY un7_0_8_cry_28(.DI(GND),.CI(un7_0_8_cry_27),.S(un7_0_8_axb_28),.O(un7_0_8_0[38:38]));
  XORCY un7_0_8_s_27(.LI(un7_0_8_axb_27),.CI(un7_0_8_cry_26),.O(un7_0_8[36:36]));
  MUXCY_L un7_0_8_cry_27_cZ(.DI(GND),.CI(un7_0_8_cry_26),.S(un7_0_8_axb_27),.LO(un7_0_8_cry_27));
  XORCY un7_0_8_s_26(.LI(un7_0_8_axb_26),.CI(un7_0_8_cry_25),.O(un7_0_8[35:35]));
  MUXCY_L un7_0_8_cry_26_cZ(.DI(GND),.CI(un7_0_8_cry_25),.S(un7_0_8_axb_26),.LO(un7_0_8_cry_26));
  XORCY un7_0_8_s_25(.LI(un7_0_8_axb_25),.CI(un7_0_8_cry_24),.O(un7_0_8[34:34]));
  MUXCY_L un7_0_8_cry_25_cZ(.DI(GND),.CI(un7_0_8_cry_24),.S(un7_0_8_axb_25),.LO(un7_0_8_cry_25));
  XORCY un7_0_8_s_24(.LI(un7_0_8_axb_24),.CI(un7_0_8_cry_23),.O(un7_0_8[33:33]));
  MUXCY_L un7_0_8_cry_24_cZ(.DI(GND),.CI(un7_0_8_cry_23),.S(un7_0_8_axb_24),.LO(un7_0_8_cry_24));
  XORCY un7_0_8_s_23(.LI(un7_0_8_axb_23),.CI(un7_0_8_cry_22),.O(un7_0_8[32:32]));
  MUXCY_L un7_0_8_cry_23_cZ(.DI(GND),.CI(un7_0_8_cry_22),.S(un7_0_8_axb_23),.LO(un7_0_8_cry_23));
  XORCY un7_0_8_s_22(.LI(un7_0_8_axb_22),.CI(un7_0_8_cry_21),.O(un7_0_8[31:31]));
  MUXCY_L un7_0_8_cry_22_cZ(.DI(GND),.CI(un7_0_8_cry_21),.S(un7_0_8_axb_22),.LO(un7_0_8_cry_22));
  XORCY un7_0_8_s_21(.LI(un7_0_8_axb_21),.CI(un7_0_8_cry_20),.O(un7_0_8[30:30]));
  MUXCY_L un7_0_8_cry_21_cZ(.DI(un7_0_8_22),.CI(un7_0_8_cry_20),.S(un7_0_8_axb_21),.LO(un7_0_8_cry_21));
  XORCY un7_0_8_s_20(.LI(un7_0_8_axb_20),.CI(un7_0_8_cry_19),.O(un7_0_8[29:29]));
  MUXCY_L un7_0_8_cry_20_cZ(.DI(un7_0_8_19),.CI(un7_0_8_cry_19),.S(un7_0_8_axb_20),.LO(un7_0_8_cry_20));
  XORCY un7_0_8_s_19(.LI(un7_0_8_axb_19),.CI(un7_0_8_cry_18),.O(un7_0_8[28:28]));
  MUXCY_L un7_0_8_cry_19_cZ(.DI(un7_0_8_cry_19_RNO),.CI(un7_0_8_cry_18),.S(un7_0_8_axb_19),.LO(un7_0_8_cry_19));
  XORCY un7_0_8_s_18(.LI(un7_0_8_axb_18),.CI(un7_0_8_cry_17),.O(un7_0_8[27:27]));
  MUXCY_L un7_0_8_cry_18_cZ(.DI(un7_0_8_cry_18_RNO),.CI(un7_0_8_cry_17),.S(un7_0_8_axb_18),.LO(un7_0_8_cry_18));
  XORCY un7_0_8_s_17(.LI(un7_0_8_axb_17),.CI(un7_0_8_cry_16),.O(un7_0_8[26:26]));
  MUXCY_L un7_0_8_cry_17_cZ(.DI(un7_0_8_cry_17_RNO),.CI(un7_0_8_cry_16),.S(un7_0_8_axb_17),.LO(un7_0_8_cry_17));
  XORCY un7_0_8_s_16(.LI(un7_0_8_axb_16),.CI(un7_0_8_cry_15),.O(un7_0_8[25:25]));
  MUXCY_L un7_0_8_cry_16_cZ(.DI(un7_0_8_cry_16_RNO),.CI(un7_0_8_cry_15),.S(un7_0_8_axb_16),.LO(un7_0_8_cry_16));
  XORCY un7_0_8_s_15(.LI(un7_0_8_axb_15),.CI(un7_0_8_cry_14),.O(un7_0_8[24:24]));
  MUXCY_L un7_0_8_cry_15_cZ(.DI(un7_0_8_cry_15_RNO),.CI(un7_0_8_cry_14),.S(un7_0_8_axb_15),.LO(un7_0_8_cry_15));
  XORCY un7_0_8_s_14(.LI(un7_0_8_axb_14),.CI(un7_0_8_cry_13),.O(un7_0_8[23:23]));
  MUXCY_L un7_0_8_cry_14_cZ(.DI(un7_0_8_cry_14_RNO),.CI(un7_0_8_cry_13),.S(un7_0_8_axb_14),.LO(un7_0_8_cry_14));
  XORCY un7_0_8_s_13(.LI(un7_0_8_axb_13),.CI(un7_0_8_cry_12),.O(un7_0_8[22:22]));
  MUXCY_L un7_0_8_cry_13_cZ(.DI(un7_0_8_cry_13_RNO),.CI(un7_0_8_cry_12),.S(un7_0_8_axb_13),.LO(un7_0_8_cry_13));
  XORCY un7_0_8_s_12(.LI(un7_0_8_axb_12),.CI(un7_0_8_cry_11),.O(un7_0_8[21:21]));
  MUXCY_L un7_0_8_cry_12_cZ(.DI(un7_0_8_cry_12_RNO),.CI(un7_0_8_cry_11),.S(un7_0_8_axb_12),.LO(un7_0_8_cry_12));
  XORCY un7_0_8_s_11(.LI(un7_0_8_axb_11),.CI(un7_0_8_cry_10),.O(un7_0_8[20:20]));
  MUXCY_L un7_0_8_cry_11_cZ(.DI(un7_0_8_cry_11_RNO),.CI(un7_0_8_cry_10),.S(un7_0_8_axb_11),.LO(un7_0_8_cry_11));
  XORCY un7_0_8_s_10(.LI(un7_0_8_axb_10),.CI(un7_0_8_cry_9),.O(un7_0_8[19:19]));
  MUXCY_L un7_0_8_cry_10_cZ(.DI(un7_0_8_cry_10_RNO),.CI(un7_0_8_cry_9),.S(un7_0_8_axb_10),.LO(un7_0_8_cry_10));
  XORCY un7_0_8_s_9(.LI(un7_0_8_axb_9),.CI(un7_0_8_cry_8),.O(un7_0_8[18:18]));
  MUXCY_L un7_0_8_cry_9_cZ(.DI(un7_0_8_cry_9_RNO),.CI(un7_0_8_cry_8),.S(un7_0_8_axb_9),.LO(un7_0_8_cry_9));
  XORCY un7_0_8_s_8(.LI(un7_0_8_axb_8),.CI(un7_0_8_cry_7),.O(un7_0_8[17:17]));
  MUXCY_L un7_0_8_cry_8_cZ(.DI(un7_0_8_cry_8_RNO),.CI(un7_0_8_cry_7),.S(un7_0_8_axb_8),.LO(un7_0_8_cry_8));
  XORCY un7_0_8_s_7(.LI(un7_0_8_axb_7),.CI(un7_0_8_cry_6),.O(un7_0_8[16:16]));
  MUXCY_L un7_0_8_cry_7_cZ(.DI(un7_0_8_cry_7_RNO),.CI(un7_0_8_cry_6),.S(un7_0_8_axb_7),.LO(un7_0_8_cry_7));
  XORCY un7_0_8_s_6(.LI(un7_0_8_axb_6),.CI(un7_0_8_cry_5),.O(un7_0_8[15:15]));
  MUXCY_L un7_0_8_cry_6_cZ(.DI(un7_0_8_cry_6_RNO),.CI(un7_0_8_cry_5),.S(un7_0_8_axb_6),.LO(un7_0_8_cry_6));
  XORCY un7_0_8_s_5(.LI(un7_0_8_axb_5),.CI(un7_0_8_cry_4),.O(un7_0_8[14:14]));
  MUXCY_L un7_0_8_cry_5_cZ(.DI(GND),.CI(un7_0_8_cry_4),.S(un7_0_8_axb_5),.LO(un7_0_8_cry_5));
  XORCY un7_0_8_s_4(.LI(un7_0_8_axb_4),.CI(un7_0_8_cry_3),.O(un7_0_8[13:13]));
  MUXCY_L un7_0_8_cry_4_cZ(.DI(ZFF_X1_10_rep1),.CI(un7_0_8_cry_3),.S(un7_0_8_axb_4),.LO(un7_0_8_cry_4));
  XORCY un7_0_8_s_3(.LI(un7_0_8_axb_3),.CI(un7_0_8_cry_2),.O(un7_0_8[12:12]));
  MUXCY_L un7_0_8_cry_3_cZ(.DI(ZFF_X1_9_rep1),.CI(un7_0_8_cry_2),.S(un7_0_8_axb_3),.LO(un7_0_8_cry_3));
  XORCY un7_0_8_s_2(.LI(un7_0_8_axb_2),.CI(un7_0_8_cry_1),.O(un7_0_8[11:11]));
  MUXCY_L un7_0_8_cry_2_cZ(.DI(ZFF_X1_5_rep1),.CI(un7_0_8_cry_1),.S(un7_0_8_axb_2),.LO(un7_0_8_cry_2));
  XORCY un7_0_8_s_1(.LI(un7_0_8_axb_1),.CI(un7_0_8_cry_0),.O(un7_0_8[10:10]));
  MUXCY_L un7_0_8_cry_1_cZ(.DI(ZFF_X1_4_rep1),.CI(un7_0_8_cry_0),.S(un7_0_8_axb_1),.LO(un7_0_8_cry_1));
  MUXCY_L un7_0_8_cry_0_cZ(.DI(ZFF_X1_fast[0:0]),.CI(GND),.S(un7_0_8[9:9]),.LO(un7_0_8_cry_0));
  XORCY un7_0_6_s_29(.LI(un7_0_6_axb_29),.CI(un7_0_6_cry_28),.O(un7_0_6[32:32]));
  MUXCY un7_0_6_cry_29(.DI(GND),.CI(un7_0_6_cry_28),.S(un7_0_6_axb_29),.O(un7_0_6_0[33:33]));
  XORCY un7_0_6_s_28(.LI(un7_0_6_axb_28),.CI(un7_0_6_cry_27),.O(un7_0_6[31:31]));
  MUXCY_L un7_0_6_cry_28_cZ(.DI(GND),.CI(un7_0_6_cry_27),.S(un7_0_6_axb_28),.LO(un7_0_6_cry_28));
  XORCY un7_0_6_s_27(.LI(un7_0_6_axb_27),.CI(un7_0_6_cry_26),.O(un7_0_6[30:30]));
  MUXCY_L un7_0_6_cry_27_cZ(.DI(GND),.CI(un7_0_6_cry_26),.S(un7_0_6_axb_27),.LO(un7_0_6_cry_27));
  XORCY un7_0_6_s_26(.LI(un7_0_6_axb_26),.CI(un7_0_6_cry_25),.O(un7_0_6[29:29]));
  MUXCY_L un7_0_6_cry_26_cZ(.DI(GND),.CI(un7_0_6_cry_25),.S(un7_0_6_axb_26),.LO(un7_0_6_cry_26));
  XORCY un7_0_6_s_25(.LI(un7_0_6_axb_25),.CI(un7_0_6_cry_24),.O(un7_0_6[28:28]));
  MUXCY_L un7_0_6_cry_25_cZ(.DI(GND),.CI(un7_0_6_cry_24),.S(un7_0_6_axb_25),.LO(un7_0_6_cry_25));
  XORCY un7_0_6_s_24(.LI(un7_0_6_axb_24),.CI(un7_0_6_cry_23),.O(un7_0_6[27:27]));
  MUXCY_L un7_0_6_cry_24_cZ(.DI(ZFF_X1[16:16]),.CI(un7_0_6_cry_23),.S(un7_0_6_axb_24),.LO(un7_0_6_cry_24));
  XORCY un7_0_6_s_23(.LI(un7_0_6_axb_23),.CI(un7_0_6_cry_22),.O(un7_0_6[26:26]));
  MUXCY_L un7_0_6_cry_23_cZ(.DI(un7_0_6_cry_23_RNO),.CI(un7_0_6_cry_22),.S(un7_0_6_axb_23),.LO(un7_0_6_cry_23));
  XORCY un7_0_6_s_22(.LI(un7_0_6_axb_22),.CI(un7_0_6_cry_21),.O(un7_0_6[25:25]));
  MUXCY_L un7_0_6_cry_22_cZ(.DI(un7_0_6_cry_22_RNO),.CI(un7_0_6_cry_21),.S(un7_0_6_axb_22),.LO(un7_0_6_cry_22));
  XORCY un7_0_6_s_21(.LI(un7_0_6_axb_21),.CI(un7_0_6_cry_20),.O(un7_0_6[24:24]));
  MUXCY_L un7_0_6_cry_21_cZ(.DI(un7_0_6_o5_20),.CI(un7_0_6_cry_20),.S(un7_0_6_axb_21),.LO(un7_0_6_cry_21));
  XORCY un7_0_6_s_20(.LI(un7_0_6_axb_20),.CI(un7_0_6_cry_19),.O(un7_0_6[23:23]));
  MUXCY_L un7_0_6_cry_20_cZ(.DI(un7_0_6_o5_19),.CI(un7_0_6_cry_19),.S(un7_0_6_axb_20),.LO(un7_0_6_cry_20));
  XORCY un7_0_6_s_19(.LI(un7_0_6_axb_19),.CI(un7_0_6_cry_18),.O(un7_0_6[22:22]));
  MUXCY_L un7_0_6_cry_19_cZ(.DI(un7_0_6_o5_18),.CI(un7_0_6_cry_18),.S(un7_0_6_axb_19),.LO(un7_0_6_cry_19));
  XORCY un7_0_6_s_18(.LI(un7_0_6_axb_18),.CI(un7_0_6_cry_17),.O(un7_0_6[21:21]));
  MUXCY_L un7_0_6_cry_18_cZ(.DI(un7_0_6_o5_17),.CI(un7_0_6_cry_17),.S(un7_0_6_axb_18),.LO(un7_0_6_cry_18));
  XORCY un7_0_6_s_17(.LI(un7_0_6_axb_17),.CI(un7_0_6_cry_16),.O(un7_0_6[20:20]));
  MUXCY_L un7_0_6_cry_17_cZ(.DI(un7_0_6_o5_16),.CI(un7_0_6_cry_16),.S(un7_0_6_axb_17),.LO(un7_0_6_cry_17));
  XORCY un7_0_6_s_16(.LI(un7_0_6_axb_16),.CI(un7_0_6_cry_15),.O(un7_0_6[19:19]));
  MUXCY_L un7_0_6_cry_16_cZ(.DI(un7_0_6_o5_15),.CI(un7_0_6_cry_15),.S(un7_0_6_axb_16),.LO(un7_0_6_cry_16));
  XORCY un7_0_6_s_15(.LI(un7_0_6_axb_15),.CI(un7_0_6_cry_14),.O(un7_0_6[18:18]));
  MUXCY_L un7_0_6_cry_15_cZ(.DI(un7_0_6_cry_15_RNO),.CI(un7_0_6_cry_14),.S(un7_0_6_axb_15),.LO(un7_0_6_cry_15));
  XORCY un7_0_6_s_14(.LI(un7_0_6_axb_14),.CI(un7_0_6_cry_13),.O(un7_0_6[17:17]));
  MUXCY_L un7_0_6_cry_14_cZ(.DI(un7_0_6_cry_14_RNO),.CI(un7_0_6_cry_13),.S(un7_0_6_axb_14),.LO(un7_0_6_cry_14));
  XORCY un7_0_6_s_13(.LI(un7_0_6_axb_13),.CI(un7_0_6_cry_12),.O(un7_0_6[16:16]));
  MUXCY_L un7_0_6_cry_13_cZ(.DI(un7_0_6_cry_13_RNO),.CI(un7_0_6_cry_12),.S(un7_0_6_axb_13),.LO(un7_0_6_cry_13));
  XORCY un7_0_6_s_12(.LI(un7_0_6_axb_12),.CI(un7_0_6_cry_11),.O(un7_0_6[15:15]));
  MUXCY_L un7_0_6_cry_12_cZ(.DI(un7_0_6_cry_12_RNO),.CI(un7_0_6_cry_11),.S(un7_0_6_axb_12),.LO(un7_0_6_cry_12));
  XORCY un7_0_6_s_11(.LI(un7_0_6_axb_11),.CI(un7_0_6_cry_10),.O(un7_0_6[14:14]));
  MUXCY_L un7_0_6_cry_11_cZ(.DI(un7_0_6_cry_11_RNO),.CI(un7_0_6_cry_10),.S(un7_0_6_axb_11),.LO(un7_0_6_cry_11));
  XORCY un7_0_6_s_10(.LI(un7_0_6_axb_10),.CI(un7_0_6_cry_9),.O(un7_0_6[13:13]));
  MUXCY_L un7_0_6_cry_10_cZ(.DI(un7_0_6_cry_10_RNO),.CI(un7_0_6_cry_9),.S(un7_0_6_axb_10),.LO(un7_0_6_cry_10));
  XORCY un7_0_6_s_9(.LI(un7_0_6_axb_9),.CI(un7_0_6_cry_8),.O(un7_0_6[12:12]));
  MUXCY_L un7_0_6_cry_9_cZ(.DI(un7_0_6_cry_9_RNO),.CI(un7_0_6_cry_8),.S(un7_0_6_axb_9),.LO(un7_0_6_cry_9));
  XORCY un7_0_6_s_8(.LI(un7_0_6_axb_8),.CI(un7_0_6_cry_7),.O(un7_0_6[11:11]));
  MUXCY_L un7_0_6_cry_8_cZ(.DI(un7_0_6_cry_8_RNO),.CI(un7_0_6_cry_7),.S(un7_0_6_axb_8),.LO(un7_0_6_cry_8));
  XORCY un7_0_6_s_7(.LI(un7_0_6_axb_7),.CI(un7_0_6_cry_6),.O(un7_0_6[10:10]));
  MUXCY_L un7_0_6_cry_7_cZ(.DI(un7_0_10_14),.CI(un7_0_6_cry_6),.S(un7_0_6_axb_7),.LO(un7_0_6_cry_7));
  XORCY un7_0_6_s_6(.LI(un7_0_6_axb_6),.CI(un7_0_6_cry_5),.O(un7_0_6[9:9]));
  MUXCY_L un7_0_6_cry_6_cZ(.DI(un7_0_6_cry_6_RNO),.CI(un7_0_6_cry_5),.S(un7_0_6_axb_6),.LO(un7_0_6_cry_6));
  XORCY un7_0_6_s_5(.LI(un7_0_6_axb_5),.CI(un7_0_6_cry_4),.O(un7_0_6[8:8]));
  MUXCY_L un7_0_6_cry_5_cZ(.DI(un7_0_6_cry_5_RNO),.CI(un7_0_6_cry_4),.S(un7_0_6_axb_5),.LO(un7_0_6_cry_5));
  XORCY un7_0_6_s_4(.LI(un7_0_6_axb_4),.CI(un7_0_6_cry_3),.O(un7_0_6[7:7]));
  MUXCY_L un7_0_6_cry_4_cZ(.DI(un7_0_6_cry_4_RNO),.CI(un7_0_6_cry_3),.S(un7_0_6_axb_4),.LO(un7_0_6_cry_4));
  XORCY un7_0_6_s_3(.LI(un7_0_6_axb_3),.CI(un7_0_6_cry_2),.O(un7_0_6[6:6]));
  MUXCY_L un7_0_6_cry_3_cZ(.DI(N_3313_i),.CI(un7_0_6_cry_2),.S(un7_0_6_axb_3),.LO(un7_0_6_cry_3));
  XORCY un7_0_6_s_2(.LI(un7_0_6_axb_2),.CI(un7_0_6_cry_1),.O(un7_0_6[5:5]));
  MUXCY_L un7_0_6_cry_2_cZ(.DI(ZFF_X1_2_rep1),.CI(un7_0_6_cry_1),.S(un7_0_6_axb_2),.LO(un7_0_6_cry_2));
  XORCY un7_0_6_s_1(.LI(un7_0_6_axb_1),.CI(un7_0_6_cry_0),.O(un7_0_6[4:4]));
  MUXCY_L un7_0_6_cry_1_cZ(.DI(ZFF_X1_fast[1:1]),.CI(un7_0_6_cry_0),.S(un7_0_6_axb_1),.LO(un7_0_6_cry_1));
  MUXCY_L un7_0_6_cry_0_cZ(.DI(ZFF_X1_0_rep1),.CI(GND),.S(un7_0_6[3:3]),.LO(un7_0_6_cry_0));
  XORCY un7_0_0_s_45_cZ(.LI(un7_0_0_axb_45),.CI(un7_0_0_cry_44),.O(un7_0_0_s_45));
  XORCY un7_0_0_s_44_cZ(.LI(un7_0_0_axb_44),.CI(un7_0_0_cry_43),.O(un7_0_0_s_44));
  MUXCY_L un7_0_0_cry_44_cZ(.DI(un7_0_10[44:44]),.CI(un7_0_0_cry_43),.S(un7_0_0_axb_44),.LO(un7_0_0_cry_44));
  XORCY un7_0_0_s_43_cZ(.LI(un7_0_0_axb_43),.CI(un7_0_0_cry_42),.O(un7_0_0_s_43));
  MUXCY_L un7_0_0_cry_43_cZ(.DI(GND),.CI(un7_0_0_cry_42),.S(un7_0_0_axb_43),.LO(un7_0_0_cry_43));
  XORCY un7_0_0_s_42_cZ(.LI(un7_0_0_axb_42),.CI(un7_0_0_cry_41),.O(un7_0_0_s_42));
  MUXCY_L un7_0_0_cry_42_cZ(.DI(GND),.CI(un7_0_0_cry_41),.S(un7_0_0_axb_42),.LO(un7_0_0_cry_42));
  XORCY un7_0_0_s_41_cZ(.LI(un7_0_0_axb_41),.CI(un7_0_0_cry_40),.O(un7_0_0_s_41));
  MUXCY_L un7_0_0_cry_41_cZ(.DI(un7_0_0_cry_41_RNO),.CI(un7_0_0_cry_40),.S(un7_0_0_axb_41),.LO(un7_0_0_cry_41));
  XORCY un7_0_0_s_40_cZ(.LI(un7_0_0_axb_40),.CI(un7_0_0_cry_39),.O(un7_0_0_s_40));
  MUXCY_L un7_0_0_cry_40_cZ(.DI(un7_0_0_cry_40_RNO),.CI(un7_0_0_cry_39),.S(un7_0_0_axb_40),.LO(un7_0_0_cry_40));
  XORCY un7_0_0_s_39_cZ(.LI(un7_0_0_axb_39),.CI(un7_0_0_cry_38),.O(un7_0_0_s_39));
  MUXCY_L un7_0_0_cry_39_cZ(.DI(un7_0_0_cry_39_RNO),.CI(un7_0_0_cry_38),.S(un7_0_0_axb_39),.LO(un7_0_0_cry_39));
  XORCY un7_0_0_s_38_cZ(.LI(un7_0_0_axb_38),.CI(un7_0_0_cry_37),.O(un7_0_0_s_38));
  MUXCY_L un7_0_0_cry_38_cZ(.DI(un7_0_0_cry_38_RNO),.CI(un7_0_0_cry_37),.S(un7_0_0_axb_38),.LO(un7_0_0_cry_38));
  XORCY un7_0_0_s_37_cZ(.LI(un7_0_0_axb_37),.CI(un7_0_0_cry_36),.O(un7_0_0_s_37));
  MUXCY_L un7_0_0_cry_37_cZ(.DI(un7_0_0_cry_37_RNO),.CI(un7_0_0_cry_36),.S(un7_0_0_axb_37),.LO(un7_0_0_cry_37));
  XORCY un7_0_0_s_36_cZ(.LI(un7_0_0_axb_36),.CI(un7_0_0_cry_35),.O(un7_0_0_s_36));
  MUXCY_L un7_0_0_cry_36_cZ(.DI(un7_0_0_cry_36_RNO),.CI(un7_0_0_cry_35),.S(un7_0_0_axb_36),.LO(un7_0_0_cry_36));
  XORCY un7_0_0_s_35_cZ(.LI(un7_0_0_axb_35),.CI(un7_0_0_cry_34),.O(un7_0_0_s_35));
  MUXCY_L un7_0_0_cry_35_cZ(.DI(un7_0_0_cry_35_RNO),.CI(un7_0_0_cry_34),.S(un7_0_0_axb_35),.LO(un7_0_0_cry_35));
  XORCY un7_0_0_s_34_cZ(.LI(un7_0_0_axb_34),.CI(un7_0_0_cry_33),.O(un7_0_0_s_34));
  MUXCY_L un7_0_0_cry_34_cZ(.DI(un7_0_0_cry_34_RNO),.CI(un7_0_0_cry_33),.S(un7_0_0_axb_34),.LO(un7_0_0_cry_34));
  XORCY un7_0_0_s_33_cZ(.LI(un7_0_0_axb_33),.CI(un7_0_0_cry_32),.O(un7_0_0_s_33));
  MUXCY_L un7_0_0_cry_33_cZ(.DI(un7_0_0_o5_32),.CI(un7_0_0_cry_32),.S(un7_0_0_axb_33),.LO(un7_0_0_cry_33));
  XORCY un7_0_0_s_32_cZ(.LI(un7_0_0_axb_32),.CI(un7_0_0_cry_31),.O(un7_0_0_s_32));
  MUXCY_L un7_0_0_cry_32_cZ(.DI(un7_0_0_o5_31),.CI(un7_0_0_cry_31),.S(un7_0_0_axb_32),.LO(un7_0_0_cry_32));
  XORCY un7_0_0_s_31_cZ(.LI(un7_0_0_axb_31),.CI(un7_0_0_cry_30),.O(un7_0_0_s_31));
  MUXCY_L un7_0_0_cry_31_cZ(.DI(un7_0_0_o5_30),.CI(un7_0_0_cry_30),.S(un7_0_0_axb_31),.LO(un7_0_0_cry_31));
  XORCY un7_0_0_s_30_cZ(.LI(un7_0_0_axb_30),.CI(un7_0_0_cry_29),.O(un7_0_0_s_30));
  MUXCY_L un7_0_0_cry_30_cZ(.DI(un7_0_0_o5_29),.CI(un7_0_0_cry_29),.S(un7_0_0_axb_30),.LO(un7_0_0_cry_30));
  XORCY un7_0_0_s_29_cZ(.LI(un7_0_0_axb_29),.CI(un7_0_0_cry_28),.O(un7_0_0_s_29));
  MUXCY_L un7_0_0_cry_29_cZ(.DI(un7_0_0_o5_28),.CI(un7_0_0_cry_28),.S(un7_0_0_axb_29),.LO(un7_0_0_cry_29));
  MUXCY_L un7_0_0_cry_28_cZ(.DI(un7_0_0_o5_27),.CI(un7_0_0_cry_27),.S(un7_0_0_axb_28),.LO(un7_0_0_cry_28));
  MUXCY_L un7_0_0_cry_27_cZ(.DI(un7_0_0_o5_26),.CI(un7_0_0_cry_26),.S(un7_0_0_axb_27),.LO(un7_0_0_cry_27));
  MUXCY_L un7_0_0_cry_26_cZ(.DI(un7_0_0_o5_25),.CI(un7_0_0_cry_25),.S(un7_0_0_axb_26),.LO(un7_0_0_cry_26));
  MUXCY_L un7_0_0_cry_25_cZ(.DI(un7_0_0_o5_24),.CI(un7_0_0_cry_24),.S(un7_0_0_axb_25),.LO(un7_0_0_cry_25));
  MUXCY_L un7_0_0_cry_24_cZ(.DI(un7_0_0_o5_23),.CI(un7_0_0_cry_23),.S(un7_0_0_axb_24),.LO(un7_0_0_cry_24));
  MUXCY_L un7_0_0_cry_23_cZ(.DI(un7_0_0_o5_22),.CI(un7_0_0_cry_22),.S(un7_0_0_axb_23),.LO(un7_0_0_cry_23));
  MUXCY_L un7_0_0_cry_22_cZ(.DI(un7_0_0_o5_21),.CI(un7_0_0_cry_21),.S(un7_0_0_axb_22),.LO(un7_0_0_cry_22));
  MUXCY_L un7_0_0_cry_21_cZ(.DI(un7_0_0_o5_20),.CI(un7_0_0_cry_20),.S(un7_0_0_axb_21),.LO(un7_0_0_cry_21));
  MUXCY_L un7_0_0_cry_20_cZ(.DI(un7_0_0_o5_19),.CI(un7_0_0_cry_19),.S(un7_0_0_axb_20),.LO(un7_0_0_cry_20));
  MUXCY_L un7_0_0_cry_19_cZ(.DI(un7_0_0_o5_18),.CI(un7_0_0_cry_18),.S(un7_0_0_axb_19),.LO(un7_0_0_cry_19));
  MUXCY_L un7_0_0_cry_18_cZ(.DI(un7_0_0_o5_17),.CI(un7_0_0_cry_17),.S(un7_0_0_axb_18),.LO(un7_0_0_cry_18));
  MUXCY_L un7_0_0_cry_17_cZ(.DI(un7_0_0_o5_16),.CI(un7_0_0_cry_16),.S(un7_0_0_axb_17),.LO(un7_0_0_cry_17));
  MUXCY_L un7_0_0_cry_16_cZ(.DI(un7_0_0_o5_15),.CI(un7_0_0_cry_15),.S(un7_0_0_axb_16),.LO(un7_0_0_cry_16));
  MUXCY_L un7_0_0_cry_15_cZ(.DI(un7_0_0_o5_14),.CI(un7_0_0_cry_14),.S(un7_0_0_axb_15),.LO(un7_0_0_cry_15));
  MUXCY_L un7_0_0_cry_14_cZ(.DI(un7_0_0_o5_13),.CI(un7_0_0_cry_13),.S(un7_0_0_axb_14),.LO(un7_0_0_cry_14));
  MUXCY_L un7_0_0_cry_13_cZ(.DI(un7_0_0_o5_12),.CI(un7_0_0_cry_12),.S(un7_0_0_axb_13),.LO(un7_0_0_cry_13));
  MUXCY_L un7_0_0_cry_12_cZ(.DI(un7_0_0_o5_11),.CI(un7_0_0_cry_11),.S(un7_0_0_axb_12),.LO(un7_0_0_cry_12));
  MUXCY_L un7_0_0_cry_11_cZ(.DI(un7_0_0_axb_10_lut6_2_O5),.CI(un7_0_0_cry_10),.S(un7_0_0_axb_11),.LO(un7_0_0_cry_11));
  MUXCY_L un7_0_0_cry_10_cZ(.DI(GND),.CI(un7_0_0_cry_9),.S(un7_0_0_axb_10),.LO(un7_0_0_cry_10));
  MUXCY_L un7_0_0_cry_9_cZ(.DI(un7_0_8[9:9]),.CI(un7_0_0_cry_8),.S(un7_0_0_axb_9),.LO(un7_0_0_cry_9));
  MUXCY_L un7_0_0_cry_8_cZ(.DI(un7_0_6[8:8]),.CI(un7_0_0_cry_7),.S(un7_0_0_axb_8),.LO(un7_0_0_cry_8));
  MUXCY_L un7_0_0_cry_7_cZ(.DI(GND),.CI(un7_0_0_cry_6),.S(un7_0_0_axb_7),.LO(un7_0_0_cry_7));
  MUXCY_L un7_0_0_cry_6_cZ(.DI(GND),.CI(un7_0_0_cry_5),.S(un7_0_0_axb_6),.LO(un7_0_0_cry_6));
  MUXCY_L un7_0_0_cry_5_cZ(.DI(GND),.CI(un7_0_0_cry_4),.S(un7_0_0_axb_5),.LO(un7_0_0_cry_5));
  MUXCY_L un7_0_0_cry_4_cZ(.DI(GND),.CI(un7_0_0_cry_3),.S(un7_0_0_axb_4),.LO(un7_0_0_cry_4));
  MUXCY_L un7_0_0_cry_3_cZ(.DI(GND),.CI(un7_0_0_cry_2),.S(un7_0_0_axb_3),.LO(un7_0_0_cry_3));
  MUXCY_L un7_0_0_cry_2_cZ(.DI(GND),.CI(un7_0_0_cry_1),.S(un7_0_0_axb_2),.LO(un7_0_0_cry_2));
  MUXCY_L un7_0_0_cry_1_cZ(.DI(GND),.CI(un7_0_0_cry_0),.S(un7_0_0_axb_1),.LO(un7_0_0_cry_1));
  MUXCY_L un7_0_0_cry_0_cZ(.DI(VCC),.CI(GND),.S(N_3353_i_0),.LO(un7_0_0_cry_0));
  XORCY un8_0_6_s_22(.LI(un8_0_6_axb_22),.CI(un8_0_6_cry_21),.O(un8_0_6[27:27]));
  MUXCY un8_0_6_cry_22(.DI(GND),.CI(un8_0_6_cry_21),.S(un8_0_6_axb_22),.O(un8_0_6_0[28:28]));
  XORCY un8_0_6_s_21(.LI(un8_0_6_axb_21),.CI(un8_0_6_cry_20),.O(un8_0_6[26:26]));
  MUXCY_L un8_0_6_cry_21_cZ(.DI(un8_0_6_43),.CI(un8_0_6_cry_20),.S(un8_0_6_axb_21),.LO(un8_0_6_cry_21));
  XORCY un8_0_6_s_20(.LI(un8_0_6_axb_20),.CI(un8_0_6_cry_19),.O(un8_0_6[25:25]));
  MUXCY_L un8_0_6_cry_20_cZ(.DI(un8_0_6_cry_20_RNO),.CI(un8_0_6_cry_19),.S(un8_0_6_axb_20),.LO(un8_0_6_cry_20));
  XORCY un8_0_6_s_19(.LI(un8_0_6_axb_19),.CI(un8_0_6_cry_18),.O(un8_0_6[24:24]));
  MUXCY_L un8_0_6_cry_19_cZ(.DI(un8_0_6_cry_19_RNO),.CI(un8_0_6_cry_18),.S(un8_0_6_axb_19),.LO(un8_0_6_cry_19));
  XORCY un8_0_6_s_18(.LI(un8_0_6_axb_18),.CI(un8_0_6_cry_17),.O(un8_0_6[23:23]));
  MUXCY_L un8_0_6_cry_18_cZ(.DI(un8_0_6_cry_18_RNO),.CI(un8_0_6_cry_17),.S(un8_0_6_axb_18),.LO(un8_0_6_cry_18));
  XORCY un8_0_6_s_17(.LI(un8_0_6_axb_17),.CI(un8_0_6_cry_16),.O(un8_0_6[22:22]));
  MUXCY_L un8_0_6_cry_17_cZ(.DI(un8_0_6_cry_17_RNO),.CI(un8_0_6_cry_16),.S(un8_0_6_axb_17),.LO(un8_0_6_cry_17));
  XORCY un8_0_6_s_16(.LI(un8_0_6_axb_16),.CI(un8_0_6_cry_15),.O(un8_0_6[21:21]));
  MUXCY_L un8_0_6_cry_16_cZ(.DI(un8_0_6_cry_16_RNO),.CI(un8_0_6_cry_15),.S(un8_0_6_axb_16),.LO(un8_0_6_cry_16));
  XORCY un8_0_6_s_15(.LI(un8_0_6_axb_15),.CI(un8_0_6_cry_14),.O(un8_0_6[20:20]));
  MUXCY_L un8_0_6_cry_15_cZ(.DI(un8_0_6_cry_15_RNO),.CI(un8_0_6_cry_14),.S(un8_0_6_axb_15),.LO(un8_0_6_cry_15));
  XORCY un8_0_6_s_14(.LI(un8_0_6_axb_14),.CI(un8_0_6_cry_13),.O(un8_0_6[19:19]));
  MUXCY_L un8_0_6_cry_14_cZ(.DI(un8_0_6_cry_14_RNO),.CI(un8_0_6_cry_13),.S(un8_0_6_axb_14),.LO(un8_0_6_cry_14));
  XORCY un8_0_6_s_13(.LI(un8_0_6_axb_13),.CI(un8_0_6_cry_12),.O(un8_0_6[18:18]));
  MUXCY_L un8_0_6_cry_13_cZ(.DI(un8_0_6_cry_13_RNO),.CI(un8_0_6_cry_12),.S(un8_0_6_axb_13),.LO(un8_0_6_cry_13));
  XORCY un8_0_6_s_12(.LI(un8_0_6_axb_12),.CI(un8_0_6_cry_11),.O(un8_0_6[17:17]));
  MUXCY_L un8_0_6_cry_12_cZ(.DI(un8_0_6_cry_12_RNO),.CI(un8_0_6_cry_11),.S(un8_0_6_axb_12),.LO(un8_0_6_cry_12));
  XORCY un8_0_6_s_11(.LI(un8_0_6_axb_11),.CI(un8_0_6_cry_10),.O(un8_0_6[16:16]));
  MUXCY_L un8_0_6_cry_11_cZ(.DI(un8_0_6_cry_11_RNO),.CI(un8_0_6_cry_10),.S(un8_0_6_axb_11),.LO(un8_0_6_cry_11));
  XORCY un8_0_6_s_10(.LI(un8_0_6_axb_10),.CI(un8_0_6_cry_9),.O(un8_0_6[15:15]));
  MUXCY_L un8_0_6_cry_10_cZ(.DI(un8_0_6_cry_10_RNO),.CI(un8_0_6_cry_9),.S(un8_0_6_axb_10),.LO(un8_0_6_cry_10));
  XORCY un8_0_6_s_9(.LI(un8_0_6_axb_9),.CI(un8_0_6_cry_8),.O(un8_0_6[14:14]));
  MUXCY_L un8_0_6_cry_9_cZ(.DI(un8_0_6_cry_9_RNO),.CI(un8_0_6_cry_8),.S(un8_0_6_axb_9),.LO(un8_0_6_cry_9));
  XORCY un8_0_6_s_8(.LI(un8_0_6_axb_8),.CI(un8_0_6_cry_7),.O(un8_0_6[13:13]));
  MUXCY_L un8_0_6_cry_8_cZ(.DI(un8_0_6_cry_8_RNO),.CI(un8_0_6_cry_7),.S(un8_0_6_axb_8),.LO(un8_0_6_cry_8));
  XORCY un8_0_6_s_7(.LI(un8_0_6_axb_7),.CI(un8_0_6_cry_6),.O(un8_0_6[12:12]));
  MUXCY_L un8_0_6_cry_7_cZ(.DI(un8_0_6_cry_7_RNO),.CI(un8_0_6_cry_6),.S(un8_0_6_axb_7),.LO(un8_0_6_cry_7));
  XORCY un8_0_6_s_6(.LI(un8_0_6_axb_6),.CI(un8_0_6_cry_5),.O(un8_0_6[11:11]));
  MUXCY_L un8_0_6_cry_6_cZ(.DI(un8_0_6_cry_6_RNO),.CI(un8_0_6_cry_5),.S(un8_0_6_axb_6),.LO(un8_0_6_cry_6));
  XORCY un8_0_6_s_5(.LI(un8_0_6_axb_5),.CI(un8_0_6_cry_4),.O(un8_0_6[10:10]));
  MUXCY_L un8_0_6_cry_5_cZ(.DI(un8_0_6_cry_5_RNO),.CI(un8_0_6_cry_4),.S(un8_0_6_axb_5),.LO(un8_0_6_cry_5));
  XORCY un8_0_6_s_4(.LI(un8_0_6_axb_4),.CI(un8_0_6_cry_3),.O(un8_0_6[9:9]));
  MUXCY_L un8_0_6_cry_4_cZ(.DI(un8_0_6_cry_4_RNO),.CI(un8_0_6_cry_3),.S(un8_0_6_axb_4),.LO(un8_0_6_cry_4));
  XORCY un8_0_6_s_3(.LI(un8_0_6_axb_3),.CI(un8_0_6_cry_2),.O(un8_0_6[8:8]));
  MUXCY_L un8_0_6_cry_3_cZ(.DI(N_3186_i),.CI(un8_0_6_cry_2),.S(un8_0_6_axb_3),.LO(un8_0_6_cry_3));
  XORCY un8_0_6_s_2(.LI(un8_0_6_axb_2),.CI(un8_0_6_cry_1),.O(un8_0_6[7:7]));
  MUXCY_L un8_0_6_cry_2_cZ(.DI(ZFF_X2[0:0]),.CI(un8_0_6_cry_1),.S(un8_0_6_axb_2),.LO(un8_0_6_cry_2));
  XORCY un8_0_6_s_1(.LI(un8_0_6_axb_1),.CI(un8_0_6_cry_0),.O(un8_0_6[6:6]));
  MUXCY_L un8_0_6_cry_1_cZ(.DI(ZFF_X2[1:1]),.CI(un8_0_6_cry_0),.S(un8_0_6_axb_1),.LO(un8_0_6_cry_1));
  MUXCY_L un8_0_6_cry_0_cZ(.DI(N_3193_i),.CI(GND),.S(un8_0_6_cry_0_sf),.LO(un8_0_6_cry_0));
  XORCY un8_0_0_s_43_cZ(.LI(un8_0_0_axb_43),.CI(un8_0_0_cry_42),.O(un8_0_0_s_43));
  XORCY un8_0_0_s_42_cZ(.LI(un8_0_0_axb_42),.CI(un8_0_0_cry_41),.O(un8_0_0_s_42));
  MUXCY_L un8_0_0_cry_42_cZ(.DI(un8_0_0_o5_41),.CI(un8_0_0_cry_41),.S(un8_0_0_axb_42),.LO(un8_0_0_cry_42));
  XORCY un8_0_0_s_41_cZ(.LI(un8_0_0_axb_41),.CI(un8_0_0_cry_40),.O(un8_0_0_s_41));
  MUXCY_L un8_0_0_cry_41_cZ(.DI(GND),.CI(un8_0_0_cry_40),.S(un8_0_0_axb_41),.LO(un8_0_0_cry_41));
  XORCY un8_0_0_s_40_cZ(.LI(N_1128_i),.CI(un8_0_0_cry_39),.O(un8_0_0_s_40));
  MUXCY_L un8_0_0_cry_40_cZ(.DI(VCC),.CI(un8_0_0_cry_39),.S(N_1128_i),.LO(un8_0_0_cry_40));
  XORCY un8_0_0_s_39_cZ(.LI(un8_0_0_axb_39),.CI(un8_0_0_cry_38),.O(un8_0_0_s_39));
  MUXCY_L un8_0_0_cry_39_cZ(.DI(un8_0_8[39:39]),.CI(un8_0_0_cry_38),.S(un8_0_0_axb_39),.LO(un8_0_0_cry_39));
  XORCY un8_0_0_s_38_cZ(.LI(un8_0_0_axb_38),.CI(un8_0_0_cry_37),.O(un8_0_0_s_38));
  MUXCY_L un8_0_0_cry_38_cZ(.DI(un8_0_0_o5_37),.CI(un8_0_0_cry_37),.S(un8_0_0_axb_38),.LO(un8_0_0_cry_38));
  XORCY un8_0_0_s_37_cZ(.LI(un8_0_0_axb_37),.CI(un8_0_0_cry_36),.O(un8_0_0_s_37));
  MUXCY_L un8_0_0_cry_37_cZ(.DI(un8_0_8_s_26_RNIUCD71_O5),.CI(un8_0_0_cry_36),.S(un8_0_0_axb_37),.LO(un8_0_0_cry_37));
  XORCY un8_0_0_s_36_cZ(.LI(un8_0_0_axb_36),.CI(un8_0_0_cry_35),.O(un8_0_0_s_36));
  MUXCY_L un8_0_0_cry_36_cZ(.DI(un8_0_0_cry_36_RNO),.CI(un8_0_0_cry_35),.S(un8_0_0_axb_36),.LO(un8_0_0_cry_36));
  XORCY un8_0_0_s_35_cZ(.LI(un8_0_0_axb_35),.CI(un8_0_0_cry_34),.O(un8_0_0_s_35));
  MUXCY_L un8_0_0_cry_35_cZ(.DI(un8_0_0_cry_35_RNO),.CI(un8_0_0_cry_34),.S(un8_0_0_axb_35),.LO(un8_0_0_cry_35));
  XORCY un8_0_0_s_34_cZ(.LI(un8_0_0_axb_34),.CI(un8_0_0_cry_33),.O(un8_0_0_s_34));
  MUXCY_L un8_0_0_cry_34_cZ(.DI(un8_0_0_cry_34_RNO),.CI(un8_0_0_cry_33),.S(un8_0_0_axb_34),.LO(un8_0_0_cry_34));
  XORCY un8_0_0_s_33_cZ(.LI(un8_0_0_axb_33),.CI(un8_0_0_cry_32),.O(un8_0_0_s_33));
  MUXCY_L un8_0_0_cry_33_cZ(.DI(un8_0_0_cry_33_RNO),.CI(un8_0_0_cry_32),.S(un8_0_0_axb_33),.LO(un8_0_0_cry_33));
  XORCY un8_0_0_s_32_cZ(.LI(un8_0_0_axb_32),.CI(un8_0_0_cry_31),.O(un8_0_0_s_32));
  MUXCY_L un8_0_0_cry_32_cZ(.DI(un8_0_0_cry_32_RNO),.CI(un8_0_0_cry_31),.S(un8_0_0_axb_32),.LO(un8_0_0_cry_32));
  XORCY un8_0_0_s_31_cZ(.LI(un8_0_0_axb_31),.CI(un8_0_0_cry_30),.O(un8_0_0_s_31));
  MUXCY_L un8_0_0_cry_31_cZ(.DI(un8_0_0_cry_31_RNO),.CI(un8_0_0_cry_30),.S(un8_0_0_axb_31),.LO(un8_0_0_cry_31));
  XORCY un8_0_0_s_30_cZ(.LI(un8_0_0_axb_30),.CI(un8_0_0_cry_29),.O(un8_0_0_s_30));
  MUXCY_L un8_0_0_cry_30_cZ(.DI(un8_0_0_cry_30_RNO),.CI(un8_0_0_cry_29),.S(un8_0_0_axb_30),.LO(un8_0_0_cry_30));
  XORCY un8_0_0_s_29_cZ(.LI(un8_0_0_axb_29),.CI(un8_0_0_cry_28),.O(un8_0_0_s_29));
  MUXCY_L un8_0_0_cry_29_cZ(.DI(un8_0_0_cry_29_RNO),.CI(un8_0_0_cry_28),.S(un8_0_0_axb_29),.LO(un8_0_0_cry_29));
  XORCY un8_0_0_s_28_cZ(.LI(un8_0_0_axb_28),.CI(un8_0_0_cry_27),.O(un8_0_0_s_28));
  MUXCY_L un8_0_0_cry_28_cZ(.DI(un8_0_0_o5_27),.CI(un8_0_0_cry_27),.S(un8_0_0_axb_28),.LO(un8_0_0_cry_28));
  MUXCY_L un8_0_0_cry_27_cZ(.DI(un8_0_0_o5_26),.CI(un8_0_0_cry_26),.S(un8_0_0_axb_27),.LO(un8_0_0_cry_27));
  MUXCY_L un8_0_0_cry_26_cZ(.DI(un8_0_0_o5_25),.CI(un8_0_0_cry_25),.S(un8_0_0_axb_26),.LO(un8_0_0_cry_26));
  MUXCY_L un8_0_0_cry_25_cZ(.DI(un8_0_0_o5_24),.CI(un8_0_0_cry_24),.S(un8_0_0_axb_25),.LO(un8_0_0_cry_25));
  MUXCY_L un8_0_0_cry_24_cZ(.DI(un8_0_0_o5_23),.CI(un8_0_0_cry_23),.S(un8_0_0_axb_24),.LO(un8_0_0_cry_24));
  MUXCY_L un8_0_0_cry_23_cZ(.DI(un8_0_0_o5_22),.CI(un8_0_0_cry_22),.S(un8_0_0_axb_23),.LO(un8_0_0_cry_23));
  MUXCY_L un8_0_0_cry_22_cZ(.DI(un8_0_0_o5_21),.CI(un8_0_0_cry_21),.S(un8_0_0_axb_22),.LO(un8_0_0_cry_22));
  MUXCY_L un8_0_0_cry_21_cZ(.DI(un8_0_0_o5_20),.CI(un8_0_0_cry_20),.S(un8_0_0_axb_21),.LO(un8_0_0_cry_21));
  MUXCY_L un8_0_0_cry_20_cZ(.DI(un8_0_0_o5_19),.CI(un8_0_0_cry_19),.S(un8_0_0_axb_20),.LO(un8_0_0_cry_20));
  MUXCY_L un8_0_0_cry_19_cZ(.DI(un8_0_0_o5_18),.CI(un8_0_0_cry_18),.S(un8_0_0_axb_19),.LO(un8_0_0_cry_19));
  MUXCY_L un8_0_0_cry_18_cZ(.DI(un8_0_0_o5_17),.CI(un8_0_0_cry_17),.S(un8_0_0_axb_18),.LO(un8_0_0_cry_18));
  MUXCY_L un8_0_0_cry_17_cZ(.DI(un8_0_0_o5_16),.CI(un8_0_0_cry_16),.S(un8_0_0_axb_17),.LO(un8_0_0_cry_17));
  MUXCY_L un8_0_0_cry_16_cZ(.DI(un8_0_0_o5_15),.CI(un8_0_0_cry_15),.S(un8_0_0_axb_16),.LO(un8_0_0_cry_16));
  MUXCY_L un8_0_0_cry_15_cZ(.DI(un8_0_0_o5_14),.CI(un8_0_0_cry_14),.S(un8_0_0_axb_15),.LO(un8_0_0_cry_15));
  MUXCY_L un8_0_0_cry_14_cZ(.DI(un8_0_0_o5_13),.CI(un8_0_0_cry_13),.S(un8_0_0_axb_14),.LO(un8_0_0_cry_14));
  MUXCY_L un8_0_0_cry_13_cZ(.DI(un8_0_0_o5_12),.CI(un8_0_0_cry_12),.S(un8_0_0_axb_13),.LO(un8_0_0_cry_13));
  MUXCY_L un8_0_0_cry_12_cZ(.DI(un8_0_0_axb_11_lut6_2_O5),.CI(un8_0_0_cry_11),.S(un8_0_0_axb_12),.LO(un8_0_0_cry_12));
  MUXCY_L un8_0_0_cry_11_cZ(.DI(GND),.CI(un8_0_0_cry_10),.S(un8_0_0_axb_11),.LO(un8_0_0_cry_11));
  MUXCY_L un8_0_0_cry_10_cZ(.DI(un8_0_6[10:10]),.CI(un8_0_0_cry_9),.S(un8_0_0_axb_10),.LO(un8_0_0_cry_10));
  MUXCY_L un8_0_0_cry_9_cZ(.DI(un8_0_6[9:9]),.CI(un8_0_0_cry_8),.S(un8_0_0_axb_9),.LO(un8_0_0_cry_9));
  MUXCY_L un8_0_0_cry_8_cZ(.DI(un8_0_6[8:8]),.CI(un8_0_0_cry_7),.S(un8_0_0_axb_8),.LO(un8_0_0_cry_8));
  MUXCY_L un8_0_0_cry_7_cZ(.DI(un8_0_6[7:7]),.CI(un8_0_0_cry_6),.S(un8_0_0_axb_7),.LO(un8_0_0_cry_7));
  MUXCY_L un8_0_0_cry_6_cZ(.DI(GND),.CI(un8_0_0_cry_5),.S(un8_0_0_cry_6_sf),.LO(un8_0_0_cry_6));
  MUXCY_L un8_0_0_cry_5_cZ(.DI(GND),.CI(un8_0_0_cry_4),.S(un8_0_6[5:5]),.LO(un8_0_0_cry_5));
  MUXCY_L un8_0_0_cry_4_cZ(.DI(GND),.CI(un8_0_0_cry_3),.S(N_3195_i),.LO(un8_0_0_cry_4));
  MUXCY_L un8_0_0_cry_3_cZ(.DI(GND),.CI(un8_0_0_cry_2),.S(N_3198_i),.LO(un8_0_0_cry_3));
  MUXCY_L un8_0_0_cry_2_cZ(.DI(GND),.CI(un8_0_0_cry_1),.S(N_3201_i),.LO(un8_0_0_cry_2));
  MUXCY_L un8_0_0_cry_1_cZ(.DI(GND),.CI(un8_0_0_cry_0),.S(N_3204_i),.LO(un8_0_0_cry_1));
  MUXCY_L un8_0_0_cry_0_cZ(.DI(GND),.CI(VCC),.S(N_3207_i),.LO(un8_0_0_cry_0));
  XORCY un10_6_s_26(.LI(un10_6_axb_26),.CI(un10_6_cry_25),.O(un10_6[35:35]));
  MUXCY un10_6_cry_26(.DI(un10_8_40),.CI(un10_6_cry_25),.S(un10_6_axb_26),.O(un10_6_0[36:36]));
  XORCY un10_6_s_25(.LI(un10_6_axb_25),.CI(un10_6_cry_24),.O(un10_6[34:34]));
  MUXCY_L un10_6_cry_25_cZ(.DI(un10_8_37),.CI(un10_6_cry_24),.S(un10_6_axb_25),.LO(un10_6_cry_25));
  XORCY un10_6_s_24(.LI(un10_6_axb_24),.CI(un10_6_cry_23),.O(un10_6[33:33]));
  MUXCY_L un10_6_cry_24_cZ(.DI(un10_8_34),.CI(un10_6_cry_23),.S(un10_6_axb_24),.LO(un10_6_cry_24));
  XORCY un10_6_s_23(.LI(un10_6_axb_23),.CI(un10_6_cry_22),.O(un10_6[32:32]));
  MUXCY_L un10_6_cry_23_cZ(.DI(un10_6_cry_23_RNO),.CI(un10_6_cry_22),.S(un10_6_axb_23),.LO(un10_6_cry_23));
  XORCY un10_6_s_22(.LI(un10_6_axb_22),.CI(un10_6_cry_21),.O(un10_6[31:31]));
  MUXCY_L un10_6_cry_22_cZ(.DI(un10_6_cry_22_RNO),.CI(un10_6_cry_21),.S(un10_6_axb_22),.LO(un10_6_cry_22));
  XORCY un10_6_s_21(.LI(un10_6_axb_21),.CI(un10_6_cry_20),.O(un10_6[30:30]));
  MUXCY_L un10_6_cry_21_cZ(.DI(un10_6_cry_21_RNO),.CI(un10_6_cry_20),.S(un10_6_axb_21),.LO(un10_6_cry_21));
  XORCY un10_6_s_20(.LI(un10_6_axb_20),.CI(un10_6_cry_19),.O(un10_6[29:29]));
  MUXCY_L un10_6_cry_20_cZ(.DI(un10_6_cry_20_RNO),.CI(un10_6_cry_19),.S(un10_6_axb_20),.LO(un10_6_cry_20));
  XORCY un10_6_s_19(.LI(un10_6_axb_19),.CI(un10_6_cry_18),.O(un10_6[28:28]));
  MUXCY_L un10_6_cry_19_cZ(.DI(un10_6_cry_19_RNO),.CI(un10_6_cry_18),.S(un10_6_axb_19),.LO(un10_6_cry_19));
  XORCY un10_6_s_18(.LI(un10_6_axb_18),.CI(un10_6_cry_17),.O(un10_6[27:27]));
  MUXCY_L un10_6_cry_18_cZ(.DI(un10_6_cry_18_RNO),.CI(un10_6_cry_17),.S(un10_6_axb_18),.LO(un10_6_cry_18));
  XORCY un10_6_s_17(.LI(un10_6_axb_17),.CI(un10_6_cry_16),.O(un10_6[26:26]));
  MUXCY_L un10_6_cry_17_cZ(.DI(un10_6_cry_17_RNO),.CI(un10_6_cry_16),.S(un10_6_axb_17),.LO(un10_6_cry_17));
  XORCY un10_6_s_16(.LI(un10_6_axb_16),.CI(un10_6_cry_15),.O(un10_6[25:25]));
  MUXCY_L un10_6_cry_16_cZ(.DI(un10_6_cry_16_RNO),.CI(un10_6_cry_15),.S(un10_6_axb_16),.LO(un10_6_cry_16));
  XORCY un10_6_s_15(.LI(un10_6_axb_15),.CI(un10_6_cry_14),.O(un10_6[24:24]));
  MUXCY_L un10_6_cry_15_cZ(.DI(un10_6_cry_15_RNO),.CI(un10_6_cry_14),.S(un10_6_axb_15),.LO(un10_6_cry_15));
  XORCY un10_6_s_14(.LI(un10_6_axb_14),.CI(un10_6_cry_13),.O(un10_6[23:23]));
  MUXCY_L un10_6_cry_14_cZ(.DI(un10_6_cry_14_RNO),.CI(un10_6_cry_13),.S(un10_6_axb_14),.LO(un10_6_cry_14));
  XORCY un10_6_s_13(.LI(un10_6_axb_13),.CI(un10_6_cry_12),.O(un10_6[22:22]));
  MUXCY_L un10_6_cry_13_cZ(.DI(un10_6_cry_13_RNO),.CI(un10_6_cry_12),.S(un10_6_axb_13),.LO(un10_6_cry_13));
  XORCY un10_6_s_12(.LI(un10_6_axb_12),.CI(un10_6_cry_11),.O(un10_6[21:21]));
  MUXCY_L un10_6_cry_12_cZ(.DI(un10_6_cry_12_RNO),.CI(un10_6_cry_11),.S(un10_6_axb_12),.LO(un10_6_cry_12));
  XORCY un10_6_s_11(.LI(un10_6_axb_11),.CI(un10_6_cry_10),.O(un10_6[20:20]));
  MUXCY_L un10_6_cry_11_cZ(.DI(un10_6_cry_11_RNO),.CI(un10_6_cry_10),.S(un10_6_axb_11),.LO(un10_6_cry_11));
  XORCY un10_6_s_10(.LI(un10_6_axb_10),.CI(un10_6_cry_9),.O(un10_6[19:19]));
  MUXCY_L un10_6_cry_10_cZ(.DI(un10_6_cry_10_RNO),.CI(un10_6_cry_9),.S(un10_6_axb_10),.LO(un10_6_cry_10));
  XORCY un10_6_s_9(.LI(un10_6_axb_9),.CI(un10_6_cry_8),.O(un10_6[18:18]));
  MUXCY_L un10_6_cry_9_cZ(.DI(un10_6_cry_9_RNO),.CI(un10_6_cry_8),.S(un10_6_axb_9),.LO(un10_6_cry_9));
  XORCY un10_6_s_8(.LI(un10_6_axb_8),.CI(un10_6_cry_7),.O(un10_6[17:17]));
  MUXCY_L un10_6_cry_8_cZ(.DI(un10_6_cry_8_RNO),.CI(un10_6_cry_7),.S(un10_6_axb_8),.LO(un10_6_cry_8));
  XORCY un10_6_s_7(.LI(un10_6_axb_7),.CI(un10_6_cry_6),.O(un10_6[16:16]));
  MUXCY_L un10_6_cry_7_cZ(.DI(un10_6_cry_7_RNO),.CI(un10_6_cry_6),.S(un10_6_axb_7),.LO(un10_6_cry_7));
  XORCY un10_6_s_6(.LI(un10_6_axb_6),.CI(un10_6_cry_5),.O(un10_6[15:15]));
  MUXCY_L un10_6_cry_6_cZ(.DI(un10_6_cry_6_RNO),.CI(un10_6_cry_5),.S(un10_6_axb_6),.LO(un10_6_cry_6));
  XORCY un10_6_s_5(.LI(un10_6_axb_5),.CI(un10_6_cry_4),.O(un10_6[14:14]));
  MUXCY_L un10_6_cry_5_cZ(.DI(un10_6_cry_5_RNO),.CI(un10_6_cry_4),.S(un10_6_axb_5),.LO(un10_6_cry_5));
  XORCY un10_6_s_4(.LI(un10_6_axb_4),.CI(un10_6_cry_3),.O(un10_6[13:13]));
  MUXCY_L un10_6_cry_4_cZ(.DI(un10_6_cry_4_RNO),.CI(un10_6_cry_3),.S(un10_6_axb_4),.LO(un10_6_cry_4));
  XORCY un10_6_s_3(.LI(un10_6_axb_3),.CI(un10_6_cry_2),.O(un10_6[12:12]));
  MUXCY_L un10_6_cry_3_cZ(.DI(un10_6_cry_3_RNO),.CI(un10_6_cry_2),.S(un10_6_axb_3),.LO(un10_6_cry_3));
  XORCY un10_6_s_2(.LI(un10_6_axb_2),.CI(un10_6_cry_1),.O(un10_6[11:11]));
  MUXCY_L un10_6_cry_2_cZ(.DI(un10_6_cry_2_RNO),.CI(un10_6_cry_1),.S(un10_6_axb_2),.LO(un10_6_cry_2));
  XORCY un10_6_s_1(.LI(un10_6_axb_1),.CI(un10_6_cry_0),.O(un10_6[10:10]));
  MUXCY_L un10_6_cry_1_cZ(.DI(un10_6_cry_1_RNO),.CI(un10_6_cry_0),.S(un10_6_axb_1),.LO(un10_6_cry_1));
  MUXCY_L un10_6_cry_0_cZ(.DI(un10_6_cry_0_RNO),.CI(GND),.S(un10_6_cry_0_RNO_0),.LO(un10_6_cry_0));
  XORCY un10_s_41_cZ(.LI(un10_8_i[47:47]),.CI(un10_cry_40),.O(un10_s_41));
  XORCY un10_s_40_cZ(.LI(un10_cry_40_sf),.CI(un10_cry_39),.O(un10_s_40));
  MUXCY_L un10_cry_40_cZ(.DI(VCC),.CI(un10_cry_39),.S(un10_cry_40_sf),.LO(un10_cry_40));
  XORCY un10_s_39_cZ(.LI(un10_8_i[45:45]),.CI(un10_cry_38),.O(un10_s_39));
  MUXCY_L un10_cry_39_cZ(.DI(VCC),.CI(un10_cry_38),.S(un10_8_i[45:45]),.LO(un10_cry_39));
  XORCY un10_s_38_cZ(.LI(un10_8_i[44:44]),.CI(un10_cry_37),.O(un10_s_38));
  MUXCY_L un10_cry_38_cZ(.DI(VCC),.CI(un10_cry_37),.S(un10_8_i[44:44]),.LO(un10_cry_38));
  XORCY un10_s_37_cZ(.LI(un10_axb_37),.CI(un10_cry_36),.O(un10_s_37));
  MUXCY_L un10_cry_37_cZ(.DI(un10_8[42:42]),.CI(un10_cry_36),.S(un10_axb_37),.LO(un10_cry_37));
  XORCY un10_s_36_cZ(.LI(un10_axb_36),.CI(un10_cry_35),.O(un10_s_36));
  MUXCY_L un10_cry_36_cZ(.DI(un10_8[41:41]),.CI(un10_cry_35),.S(un10_axb_36),.LO(un10_cry_36));
  XORCY un10_s_35_cZ(.LI(un10_axb_35),.CI(un10_cry_34),.O(un10_s_35));
  MUXCY_L un10_cry_35_cZ(.DI(un10_8[40:40]),.CI(un10_cry_34),.S(un10_axb_35),.LO(un10_cry_35));
  XORCY un10_s_34_cZ(.LI(un10_axb_34),.CI(un10_cry_33),.O(un10_s_34));
  MUXCY_L un10_cry_34_cZ(.DI(un10_8[39:39]),.CI(un10_cry_33),.S(un10_axb_34),.LO(un10_cry_34));
  XORCY un10_s_33_cZ(.LI(un10_axb_33),.CI(un10_cry_32),.O(un10_s_33));
  MUXCY_L un10_cry_33_cZ(.DI(un10_8[38:38]),.CI(un10_cry_32),.S(un10_axb_33),.LO(un10_cry_33));
  XORCY un10_s_32_cZ(.LI(un10_axb_32),.CI(un10_cry_31),.O(un10_s_32));
  MUXCY_L un10_cry_32_cZ(.DI(un10_8[37:37]),.CI(un10_cry_31),.S(un10_axb_32),.LO(un10_cry_32));
  XORCY un10_s_31_cZ(.LI(un10_axb_31),.CI(un10_cry_30),.O(un10_s_31));
  MUXCY_L un10_cry_31_cZ(.DI(un10_cry_31_RNO),.CI(un10_cry_30),.S(un10_axb_31),.LO(un10_cry_31));
  XORCY un10_s_30_cZ(.LI(un10_axb_30),.CI(un10_cry_29),.O(un10_s_30));
  MUXCY_L un10_cry_30_cZ(.DI(un10_cry_30_RNO),.CI(un10_cry_29),.S(un10_axb_30),.LO(un10_cry_30));
  XORCY un10_s_29_cZ(.LI(un10_axb_29),.CI(un10_cry_28),.O(un10_s_29));
  MUXCY_L un10_cry_29_cZ(.DI(un10_cry_29_RNO),.CI(un10_cry_28),.S(un10_axb_29),.LO(un10_cry_29));
  XORCY un10_s_28_cZ(.LI(un10_axb_28),.CI(un10_cry_27),.O(un10_s_28));
  MUXCY_L un10_cry_28_cZ(.DI(un10_o5_27),.CI(un10_cry_27),.S(un10_axb_28),.LO(un10_cry_28));
  XORCY un10_s_27_cZ(.LI(un10_axb_27),.CI(un10_cry_26),.O(un10_s_27));
  MUXCY_L un10_cry_27_cZ(.DI(un10_o5_26),.CI(un10_cry_26),.S(un10_axb_27),.LO(un10_cry_27));
  XORCY un10_s_26_cZ(.LI(un10_axb_26),.CI(un10_cry_25),.O(un10_s_26));
  MUXCY_L un10_cry_26_cZ(.DI(un10_o5_25),.CI(un10_cry_25),.S(un10_axb_26),.LO(un10_cry_26));
  XORCY un10_s_25_cZ(.LI(un10_axb_25),.CI(un10_cry_24),.O(un10_s_25));
  MUXCY_L un10_cry_25_cZ(.DI(un10_o5_24),.CI(un10_cry_24),.S(un10_axb_25),.LO(un10_cry_25));
  XORCY un10_s_24_cZ(.LI(un10_axb_24),.CI(un10_cry_23),.O(un10_s_24));
  MUXCY_L un10_cry_24_cZ(.DI(un10_o5_23),.CI(un10_cry_23),.S(un10_axb_24),.LO(un10_cry_24));
  MUXCY_L un10_cry_23_cZ(.DI(un10_o5_22),.CI(un10_cry_22),.S(un10_axb_23),.LO(un10_cry_23));
  MUXCY_L un10_cry_22_cZ(.DI(un10_o5_21),.CI(un10_cry_21),.S(un10_axb_22),.LO(un10_cry_22));
  MUXCY_L un10_cry_21_cZ(.DI(un10_o5_20),.CI(un10_cry_20),.S(un10_axb_21),.LO(un10_cry_21));
  MUXCY_L un10_cry_20_cZ(.DI(un10_o5_19),.CI(un10_cry_19),.S(un10_axb_20),.LO(un10_cry_20));
  MUXCY_L un10_cry_19_cZ(.DI(un10_o5_18),.CI(un10_cry_18),.S(un10_axb_19),.LO(un10_cry_19));
  MUXCY_L un10_cry_18_cZ(.DI(un10_o5_17),.CI(un10_cry_17),.S(un10_axb_18),.LO(un10_cry_18));
  MUXCY_L un10_cry_17_cZ(.DI(un10_o5_16),.CI(un10_cry_16),.S(un10_axb_17),.LO(un10_cry_17));
  MUXCY_L un10_cry_16_cZ(.DI(un10_o5_15),.CI(un10_cry_15),.S(un10_axb_16),.LO(un10_cry_16));
  MUXCY_L un10_cry_15_cZ(.DI(un10_o5_14),.CI(un10_cry_14),.S(un10_axb_15),.LO(un10_cry_15));
  MUXCY_L un10_cry_14_cZ(.DI(un10_o5_13),.CI(un10_cry_13),.S(un10_axb_14),.LO(un10_cry_14));
  MUXCY_L un10_cry_13_cZ(.DI(un10_o5_12),.CI(un10_cry_12),.S(un10_axb_13),.LO(un10_cry_13));
  MUXCY_L un10_cry_12_cZ(.DI(un10_axb_11_lut6_2_O5),.CI(un10_cry_11),.S(un10_axb_12),.LO(un10_cry_12));
  MUXCY_L un10_cry_11_cZ(.DI(un10_6[17:17]),.CI(un10_cry_10),.S(un10_axb_11),.LO(un10_cry_11));
  MUXCY_L un10_cry_10_cZ(.DI(un10_6[16:16]),.CI(un10_cry_9),.S(un10_axb_10),.LO(un10_cry_10));
  MUXCY_L un10_cry_9_cZ(.DI(un10_6[15:15]),.CI(un10_cry_8),.S(un10_axb_9),.LO(un10_cry_9));
  MUXCY_L un10_cry_8_cZ(.DI(un10_6[14:14]),.CI(un10_cry_7),.S(un10_axb_8),.LO(un10_cry_8));
  MUXCY_L un10_cry_7_cZ(.DI(un10_6[13:13]),.CI(un10_cry_6),.S(un10_axb_7),.LO(un10_cry_7));
  MUXCY_L un10_cry_6_cZ(.DI(un10_6[12:12]),.CI(un10_cry_5),.S(un10_axb_6),.LO(un10_cry_6));
  MUXCY_L un10_cry_5_cZ(.DI(un10_6[11:11]),.CI(un10_cry_4),.S(un10_axb_5),.LO(un10_cry_5));
  MUXCY_L un10_cry_4_cZ(.DI(un10_6[10:10]),.CI(un10_cry_3),.S(un10_axb_4),.LO(un10_cry_4));
  MUXCY_L un10_cry_3_cZ(.DI(un10_6[9:9]),.CI(un10_cry_2),.S(un10_axb_3),.LO(un10_cry_3));
  MUXCY_L un10_cry_2_cZ(.DI(un10_6[8:8]),.CI(un10_cry_1),.S(un10_axb_2),.LO(un10_cry_2));
  MUXCY_L un10_cry_1_cZ(.DI(un10_6[7:7]),.CI(un10_cry_0),.S(un10_axb_1),.LO(un10_cry_1));
  MUXCY_L un10_cry_0_cZ(.DI(un10_6[6:6]),.CI(GND),.S(un10_6_i[6:6]),.LO(un10_cry_0));
  XORCY un9_10_s_29(.LI(un9_10_axb_29),.CI(un9_10_cry_28),.O(un9_10[41:41]));
  MUXCY un9_10_cry_29(.DI(GND),.CI(un9_10_cry_28),.S(un9_10_axb_29),.O(un9_10_0[42:42]));
  XORCY un9_10_s_28(.LI(un9_10_axb_28),.CI(un9_10_cry_27),.O(un9_10[40:40]));
  MUXCY_L un9_10_cry_28_cZ(.DI(GND),.CI(un9_10_cry_27),.S(un9_10_axb_28),.LO(un9_10_cry_28));
  XORCY un9_10_s_27(.LI(un9_10_axb_27),.CI(un9_10_cry_26),.O(un9_10[39:39]));
  MUXCY_L un9_10_cry_27_cZ(.DI(un9_10_cry_27_RNO),.CI(un9_10_cry_26),.S(un9_10_axb_27),.LO(un9_10_cry_27));
  XORCY un9_10_s_26(.LI(un9_10_axb_26),.CI(un9_10_cry_25),.O(un9_10[38:38]));
  MUXCY_L un9_10_cry_26_cZ(.DI(un9_10_cry_26_RNO),.CI(un9_10_cry_25),.S(un9_10_axb_26),.LO(un9_10_cry_26));
  XORCY un9_10_s_25(.LI(un9_10_axb_25),.CI(un9_10_cry_24),.O(un9_10[37:37]));
  MUXCY_L un9_10_cry_25_cZ(.DI(un9_10_cry_25_RNO),.CI(un9_10_cry_24),.S(un9_10_axb_25),.LO(un9_10_cry_25));
  XORCY un9_10_s_24(.LI(un9_10_axb_24),.CI(un9_10_cry_23),.O(un9_10[36:36]));
  MUXCY_L un9_10_cry_24_cZ(.DI(un9_10_cry_24_RNO),.CI(un9_10_cry_23),.S(un9_10_axb_24),.LO(un9_10_cry_24));
  XORCY un9_10_s_23(.LI(un9_10_axb_23),.CI(un9_10_cry_22),.O(un9_10[35:35]));
  MUXCY_L un9_10_cry_23_cZ(.DI(un9_10_cry_23_RNO),.CI(un9_10_cry_22),.S(un9_10_axb_23),.LO(un9_10_cry_23));
  XORCY un9_10_s_22(.LI(un9_10_axb_22),.CI(un9_10_cry_21),.O(un9_10[34:34]));
  MUXCY_L un9_10_cry_22_cZ(.DI(un9_10_cry_22_RNO),.CI(un9_10_cry_21),.S(un9_10_axb_22),.LO(un9_10_cry_22));
  XORCY un9_10_s_21(.LI(un9_10_axb_21),.CI(un9_10_cry_20),.O(un9_10[33:33]));
  MUXCY_L un9_10_cry_21_cZ(.DI(un9_10_cry_21_RNO),.CI(un9_10_cry_20),.S(un9_10_axb_21),.LO(un9_10_cry_21));
  XORCY un9_10_s_20(.LI(un9_10_axb_20),.CI(un9_10_cry_19),.O(un9_10[32:32]));
  MUXCY_L un9_10_cry_20_cZ(.DI(un9_10_cry_20_RNO),.CI(un9_10_cry_19),.S(un9_10_axb_20),.LO(un9_10_cry_20));
  XORCY un9_10_s_19(.LI(un9_10_axb_19),.CI(un9_10_cry_18),.O(un9_10[31:31]));
  MUXCY_L un9_10_cry_19_cZ(.DI(un9_10_cry_19_RNO),.CI(un9_10_cry_18),.S(un9_10_axb_19),.LO(un9_10_cry_19));
  XORCY un9_10_s_18(.LI(un9_10_axb_18),.CI(un9_10_cry_17),.O(un9_10[30:30]));
  MUXCY_L un9_10_cry_18_cZ(.DI(un9_10_cry_18_RNO),.CI(un9_10_cry_17),.S(un9_10_axb_18),.LO(un9_10_cry_18));
  XORCY un9_10_s_17(.LI(un9_10_axb_17),.CI(un9_10_cry_16),.O(un9_10[29:29]));
  MUXCY_L un9_10_cry_17_cZ(.DI(un9_10_cry_17_RNO),.CI(un9_10_cry_16),.S(un9_10_axb_17),.LO(un9_10_cry_17));
  XORCY un9_10_s_16(.LI(un9_10_axb_16),.CI(un9_10_cry_15),.O(un9_10[28:28]));
  MUXCY_L un9_10_cry_16_cZ(.DI(un9_10_cry_16_RNO),.CI(un9_10_cry_15),.S(un9_10_axb_16),.LO(un9_10_cry_16));
  XORCY un9_10_s_15(.LI(un9_10_axb_15),.CI(un9_10_cry_14),.O(un9_10[27:27]));
  MUXCY_L un9_10_cry_15_cZ(.DI(un9_10_cry_15_RNO),.CI(un9_10_cry_14),.S(un9_10_axb_15),.LO(un9_10_cry_15));
  XORCY un9_10_s_14(.LI(un9_10_axb_14),.CI(un9_10_cry_13),.O(un9_10[26:26]));
  MUXCY_L un9_10_cry_14_cZ(.DI(un9_10_cry_14_RNO),.CI(un9_10_cry_13),.S(un9_10_axb_14),.LO(un9_10_cry_14));
  XORCY un9_10_s_13(.LI(un9_10_axb_13),.CI(un9_10_cry_12),.O(un9_10[25:25]));
  MUXCY_L un9_10_cry_13_cZ(.DI(un9_10_cry_13_RNO),.CI(un9_10_cry_12),.S(un9_10_axb_13),.LO(un9_10_cry_13));
  XORCY un9_10_s_12(.LI(un9_10_axb_12),.CI(un9_10_cry_11),.O(un9_10[24:24]));
  MUXCY_L un9_10_cry_12_cZ(.DI(un9_10_cry_12_RNO),.CI(un9_10_cry_11),.S(un9_10_axb_12),.LO(un9_10_cry_12));
  XORCY un9_10_s_11(.LI(un9_10_axb_11),.CI(un9_10_cry_10),.O(un9_10[23:23]));
  MUXCY_L un9_10_cry_11_cZ(.DI(un9_10_cry_11_RNO),.CI(un9_10_cry_10),.S(un9_10_axb_11),.LO(un9_10_cry_11));
  XORCY un9_10_s_10(.LI(un9_10_axb_10),.CI(un9_10_cry_9),.O(un9_10[22:22]));
  MUXCY_L un9_10_cry_10_cZ(.DI(un9_10_cry_10_RNO),.CI(un9_10_cry_9),.S(un9_10_axb_10),.LO(un9_10_cry_10));
  XORCY un9_10_s_9(.LI(un9_10_axb_9),.CI(un9_10_cry_8),.O(un9_10[21:21]));
  MUXCY_L un9_10_cry_9_cZ(.DI(un9_10_cry_9_RNO),.CI(un9_10_cry_8),.S(un9_10_axb_9),.LO(un9_10_cry_9));
  XORCY un9_10_s_8(.LI(un9_10_axb_8),.CI(un9_10_cry_7),.O(un9_10[20:20]));
  MUXCY_L un9_10_cry_8_cZ(.DI(un9_10_cry_8_RNO),.CI(un9_10_cry_7),.S(un9_10_axb_8),.LO(un9_10_cry_8));
  XORCY un9_10_s_7(.LI(un9_10_axb_7),.CI(un9_10_cry_6),.O(un9_10[19:19]));
  MUXCY_L un9_10_cry_7_cZ(.DI(un9_10_cry_7_RNO),.CI(un9_10_cry_6),.S(un9_10_axb_7),.LO(un9_10_cry_7));
  XORCY un9_10_s_6(.LI(un9_10_axb_6),.CI(un9_10_cry_5),.O(un9_10[18:18]));
  MUXCY_L un9_10_cry_6_cZ(.DI(un9_10_cry_6_RNO),.CI(un9_10_cry_5),.S(un9_10_axb_6),.LO(un9_10_cry_6));
  XORCY un9_10_s_5(.LI(un9_10_axb_5),.CI(un9_10_cry_4),.O(un9_10[17:17]));
  MUXCY_L un9_10_cry_5_cZ(.DI(un9_10_cry_5_RNO),.CI(un9_10_cry_4),.S(un9_10_axb_5),.LO(un9_10_cry_5));
  XORCY un9_10_s_4(.LI(un9_10_axb_4),.CI(un9_10_cry_3),.O(un9_10[16:16]));
  MUXCY_L un9_10_cry_4_cZ(.DI(un9_10_cry_4_RNO),.CI(un9_10_cry_3),.S(un9_10_axb_4),.LO(un9_10_cry_4));
  XORCY un9_10_s_3(.LI(un9_10_axb_3),.CI(un9_10_cry_2),.O(un9_10[15:15]));
  MUXCY_L un9_10_cry_3_cZ(.DI(un9_10_cry_3_RNO),.CI(un9_10_cry_2),.S(un9_10_axb_3),.LO(un9_10_cry_3));
  XORCY un9_10_s_2(.LI(un9_10_axb_2),.CI(un9_10_cry_1),.O(un9_10[14:14]));
  MUXCY_L un9_10_cry_2_cZ(.DI(GND),.CI(un9_10_cry_1),.S(un9_10_axb_2),.LO(un9_10_cry_2));
  XORCY un9_10_s_1(.LI(un9_10_axb_1),.CI(un9_10_cry_0),.O(un9_10[13:13]));
  MUXCY_L un9_10_cry_1_cZ(.DI(GND),.CI(un9_10_cry_0),.S(un9_10_axb_1),.LO(un9_10_cry_1));
  MUXCY_L un9_10_cry_0_cZ(.DI(un9_10_fast[8:8]),.CI(GND),.S(un9_10[12:12]),.LO(un9_10_cry_0));
  XORCY un9_8_s_35(.LI(un9_8_axb_35),.CI(un9_8_cry_34),.O(un9_8[43:43]));
  MUXCY_L un9_8_cry_35(.DI(GND),.CI(un9_8_cry_34),.S(un9_8_axb_35),.LO(un9_8[45:45]));
  XORCY un9_8_s_34(.LI(un9_8_axb_34),.CI(un9_8_cry_33),.O(un9_8[42:42]));
  MUXCY_L un9_8_cry_34_cZ(.DI(GND),.CI(un9_8_cry_33),.S(un9_8_axb_34),.LO(un9_8_cry_34));
  XORCY un9_8_s_33(.LI(un9_8_axb_33),.CI(un9_8_cry_32),.O(un9_8[41:41]));
  MUXCY_L un9_8_cry_33_cZ(.DI(GND),.CI(un9_8_cry_32),.S(un9_8_axb_33),.LO(un9_8_cry_33));
  XORCY un9_8_s_32(.LI(un9_8_axb_32),.CI(un9_8_cry_31),.O(un9_8[40:40]));
  MUXCY_L un9_8_cry_32_cZ(.DI(GND),.CI(un9_8_cry_31),.S(un9_8_axb_32),.LO(un9_8_cry_32));
  XORCY un9_8_s_31(.LI(un9_8_axb_31),.CI(un9_8_cry_30),.O(un9_8[39:39]));
  MUXCY_L un9_8_cry_31_cZ(.DI(GND),.CI(un9_8_cry_30),.S(un9_8_axb_31),.LO(un9_8_cry_31));
  MUXCY_L un9_8_cry_30_cZ(.DI(VCC),.CI(un9_8_cry_29),.S(un9_8_cry_30_RNO),.LO(un9_8_cry_30));
  XORCY un9_8_s_29(.LI(un9_8_axb_29),.CI(un9_8_cry_28),.O(un9_8[37:37]));
  XORCY un9_8_s_28(.LI(un9_8_axb_28),.CI(un9_8_cry_27),.O(un9_8[36:36]));
  MUXCY_L un9_8_cry_28_cZ(.DI(un9_11[26:26]),.CI(un9_8_cry_27),.S(un9_8_axb_28),.LO(un9_8_cry_28));
  XORCY un9_8_s_27(.LI(un9_8_axb_27),.CI(un9_8_cry_26),.O(un9_8[35:35]));
  MUXCY_L un9_8_cry_27_cZ(.DI(un9_11[25:25]),.CI(un9_8_cry_26),.S(un9_8_axb_27),.LO(un9_8_cry_27));
  XORCY un9_8_s_26(.LI(un9_8_axb_26),.CI(un9_8_cry_25),.O(un9_8[34:34]));
  MUXCY_L un9_8_cry_26_cZ(.DI(un9_11[24:24]),.CI(un9_8_cry_25),.S(un9_8_axb_26),.LO(un9_8_cry_26));
  XORCY un9_8_s_25(.LI(un9_8_axb_25),.CI(un9_8_cry_24),.O(un9_8[33:33]));
  MUXCY_L un9_8_cry_25_cZ(.DI(un9_11[23:23]),.CI(un9_8_cry_24),.S(un9_8_axb_25),.LO(un9_8_cry_25));
  XORCY un9_8_s_24(.LI(un9_8_axb_24),.CI(un9_8_cry_23),.O(un9_8[32:32]));
  MUXCY_L un9_8_cry_24_cZ(.DI(un9_11[22:22]),.CI(un9_8_cry_23),.S(un9_8_axb_24),.LO(un9_8_cry_24));
  XORCY un9_8_s_23(.LI(un9_8_axb_23),.CI(un9_8_cry_22),.O(un9_8[31:31]));
  MUXCY_L un9_8_cry_23_cZ(.DI(un9_8_cry_23_RNO),.CI(un9_8_cry_22),.S(un9_8_axb_23),.LO(un9_8_cry_23));
  XORCY un9_8_s_22(.LI(un9_8_axb_22),.CI(un9_8_cry_21),.O(un9_8[30:30]));
  MUXCY_L un9_8_cry_22_cZ(.DI(un9_8_cry_22_RNO),.CI(un9_8_cry_21),.S(un9_8_axb_22),.LO(un9_8_cry_22));
  XORCY un9_8_s_21(.LI(un9_8_axb_21),.CI(un9_8_cry_20),.O(un9_8[29:29]));
  MUXCY_L un9_8_cry_21_cZ(.DI(un9_8_cry_21_RNO),.CI(un9_8_cry_20),.S(un9_8_axb_21),.LO(un9_8_cry_21));
  XORCY un9_8_s_20(.LI(un9_8_axb_20),.CI(un9_8_cry_19),.O(un9_8[28:28]));
  MUXCY_L un9_8_cry_20_cZ(.DI(un9_8_o5_19),.CI(un9_8_cry_19),.S(un9_8_axb_20),.LO(un9_8_cry_20));
  XORCY un9_8_s_19(.LI(un9_8_axb_19),.CI(un9_8_cry_18),.O(un9_8[27:27]));
  MUXCY_L un9_8_cry_19_cZ(.DI(un9_8_o5_18),.CI(un9_8_cry_18),.S(un9_8_axb_19),.LO(un9_8_cry_19));
  XORCY un9_8_s_18(.LI(un9_8_axb_18),.CI(un9_8_cry_17),.O(un9_8[26:26]));
  MUXCY_L un9_8_cry_18_cZ(.DI(un9_8_o5_17),.CI(un9_8_cry_17),.S(un9_8_axb_18),.LO(un9_8_cry_18));
  XORCY un9_8_s_17(.LI(un9_8_axb_17),.CI(un9_8_cry_16),.O(un9_8[25:25]));
  MUXCY_L un9_8_cry_17_cZ(.DI(un9_8_cry_17_RNO),.CI(un9_8_cry_16),.S(un9_8_axb_17),.LO(un9_8_cry_17));
  XORCY un9_8_s_16(.LI(un9_8_axb_16),.CI(un9_8_cry_15),.O(un9_8[24:24]));
  MUXCY_L un9_8_cry_16_cZ(.DI(un9_8_o5_15),.CI(un9_8_cry_15),.S(un9_8_axb_16),.LO(un9_8_cry_16));
  XORCY un9_8_s_15(.LI(un9_8_axb_15),.CI(un9_8_cry_14),.O(un9_8[23:23]));
  MUXCY_L un9_8_cry_15_cZ(.DI(un9_8_o5_14),.CI(un9_8_cry_14),.S(un9_8_axb_15),.LO(un9_8_cry_15));
  XORCY un9_8_s_14(.LI(un9_8_axb_14),.CI(un9_8_cry_13),.O(un9_8[22:22]));
  MUXCY_L un9_8_cry_14_cZ(.DI(un9_8_o5_13),.CI(un9_8_cry_13),.S(un9_8_axb_14),.LO(un9_8_cry_14));
  XORCY un9_8_s_13(.LI(un9_8_axb_13),.CI(un9_8_cry_12),.O(un9_8[21:21]));
  MUXCY_L un9_8_cry_13_cZ(.DI(un9_8_cry_13_RNO),.CI(un9_8_cry_12),.S(un9_8_axb_13),.LO(un9_8_cry_13));
  XORCY un9_8_s_12(.LI(un9_8_axb_12),.CI(un9_8_cry_11),.O(un9_8[20:20]));
  MUXCY_L un9_8_cry_12_cZ(.DI(un9_8_cry_12_RNO),.CI(un9_8_cry_11),.S(un9_8_axb_12),.LO(un9_8_cry_12));
  XORCY un9_8_s_11(.LI(un9_8_axb_11),.CI(un9_8_cry_10),.O(un9_8[19:19]));
  MUXCY_L un9_8_cry_11_cZ(.DI(un9_8_cry_11_RNO),.CI(un9_8_cry_10),.S(un9_8_axb_11),.LO(un9_8_cry_11));
  XORCY un9_8_s_10(.LI(un9_8_axb_10),.CI(un9_8_cry_9),.O(un9_8[18:18]));
  MUXCY_L un9_8_cry_10_cZ(.DI(un9_8_cry_10_RNO),.CI(un9_8_cry_9),.S(un9_8_axb_10),.LO(un9_8_cry_10));
  XORCY un9_8_s_9(.LI(un9_8_axb_9),.CI(un9_8_cry_8),.O(un9_8[17:17]));
  MUXCY_L un9_8_cry_9_cZ(.DI(un9_8_cry_9_RNO),.CI(un9_8_cry_8),.S(un9_8_axb_9),.LO(un9_8_cry_9));
  XORCY un9_8_s_8(.LI(un9_8_axb_8),.CI(un9_8_cry_7),.O(un9_8[16:16]));
  MUXCY_L un9_8_cry_8_cZ(.DI(un9_8_cry_8_RNO),.CI(un9_8_cry_7),.S(un9_8_axb_8),.LO(un9_8_cry_8));
  XORCY un9_8_s_7(.LI(un9_8_axb_7),.CI(un9_8_cry_6),.O(un9_8[15:15]));
  MUXCY_L un9_8_cry_7_cZ(.DI(un9_8_cry_7_RNO),.CI(un9_8_cry_6),.S(un9_8_axb_7),.LO(un9_8_cry_7));
  XORCY un9_8_s_6(.LI(un9_8_axb_6),.CI(un9_8_cry_5),.O(un9_8[14:14]));
  MUXCY_L un9_8_cry_6_cZ(.DI(un9_8_cry_6_RNO),.CI(un9_8_cry_5),.S(un9_8_axb_6),.LO(un9_8_cry_6));
  XORCY un9_8_s_5(.LI(un9_8_axb_5),.CI(un9_8_cry_4),.O(un9_8[13:13]));
  MUXCY_L un9_8_cry_5_cZ(.DI(un9_11_i[23:23]),.CI(un9_8_cry_4),.S(un9_8_axb_5),.LO(un9_8_cry_5));
  XORCY un9_8_s_4(.LI(un9_8_axb_4),.CI(un9_8_cry_3),.O(un9_8[12:12]));
  MUXCY_L un9_8_cry_4_cZ(.DI(ZFF_Y1_7_rep1),.CI(un9_8_cry_3),.S(un9_8_axb_4),.LO(un9_8_cry_4));
  XORCY un9_8_s_3(.LI(un9_8_axb_3),.CI(un9_8_cry_2),.O(un9_8[11:11]));
  MUXCY_L un9_8_cry_3_cZ(.DI(ZFF_Y1_3_rep1),.CI(un9_8_cry_2),.S(un9_8_axb_3),.LO(un9_8_cry_3));
  XORCY un9_8_s_2(.LI(un9_8_axb_2),.CI(un9_8_cry_1),.O(un9_8[10:10]));
  MUXCY_L un9_8_cry_2_cZ(.DI(un9_8_7_rep1),.CI(un9_8_cry_1),.S(un9_8_axb_2),.LO(un9_8_cry_2));
  XORCY un9_8_s_1(.LI(un9_8_axb_1),.CI(un9_8_cry_0),.O(un9_8[9:9]));
  MUXCY_L un9_8_cry_1_cZ(.DI(ZFF_Y1_4_rep1),.CI(un9_8_cry_0),.S(un9_8_axb_1),.LO(un9_8_cry_1));
  MUXCY_L un9_8_cry_0_cZ(.DI(ZFF_Y1_3_rep1),.CI(GND),.S(un9_8_cry_0_RNO),.LO(un9_8_cry_0));
  XORCY un9_6_0_s_46(.LI(un9_6_0_axb_46),.CI(un9_6_0_cry_45),.O(un9_6[46:46]));
  MUXCY un9_6_0_cry_46(.DI(GND),.CI(un9_6_0_cry_45),.S(un9_6_0_axb_46),.O(un9_6_0[47:47]));
  XORCY un9_6_0_s_45(.LI(un9_6_0_axb_45),.CI(un9_6_0_cry_44),.O(un9_6[45:45]));
  MUXCY_L un9_6_0_cry_45_cZ(.DI(un9_11[45:45]),.CI(un9_6_0_cry_44),.S(un9_6_0_axb_45),.LO(un9_6_0_cry_45));
  XORCY un9_6_0_s_44(.LI(un9_6_0_axb_44),.CI(un9_6_0_cry_43),.O(un9_6[44:44]));
  MUXCY_L un9_6_0_cry_44_cZ(.DI(GND),.CI(un9_6_0_cry_43),.S(un9_6_0_axb_44),.LO(un9_6_0_cry_44));
  XORCY un9_6_0_s_43(.LI(un9_6_0_axb_43),.CI(un9_6_0_cry_42),.O(un9_6[43:43]));
  MUXCY_L un9_6_0_cry_43_cZ(.DI(un9_11[43:43]),.CI(un9_6_0_cry_42),.S(un9_6_0_axb_43),.LO(un9_6_0_cry_43));
  XORCY un9_6_0_s_42(.LI(un9_6_0_axb_42),.CI(un9_6_0_cry_41),.O(un9_6[42:42]));
  MUXCY_L un9_6_0_cry_42_cZ(.DI(GND),.CI(un9_6_0_cry_41),.S(un9_6_0_axb_42),.LO(un9_6_0_cry_42));
  XORCY un9_6_0_s_41(.LI(un9_6_0_axb_41),.CI(un9_6_0_cry_40),.O(un9_6[41:41]));
  MUXCY_L un9_6_0_cry_41_cZ(.DI(un9_11[41:41]),.CI(un9_6_0_cry_40),.S(un9_6_0_axb_41),.LO(un9_6_0_cry_41));
  XORCY un9_6_0_s_40(.LI(un9_6_0_axb_40),.CI(un9_6_0_cry_39),.O(un9_6[40:40]));
  MUXCY_L un9_6_0_cry_40_cZ(.DI(un9_11[40:40]),.CI(un9_6_0_cry_39),.S(un9_6_0_axb_40),.LO(un9_6_0_cry_40));
  XORCY un9_6_0_s_39(.LI(un9_6_0_axb_39),.CI(un9_6_0_cry_38),.O(un9_6[39:39]));
  MUXCY_L un9_6_0_cry_39_cZ(.DI(GND),.CI(un9_6_0_cry_38),.S(un9_6_0_axb_39),.LO(un9_6_0_cry_39));
  XORCY un9_6_0_s_38(.LI(un9_6_0_axb_38),.CI(un9_6_0_cry_37),.O(un9_6[38:38]));
  MUXCY_L un9_6_0_cry_38_cZ(.DI(GND),.CI(un9_6_0_cry_37),.S(un9_6_0_axb_38),.LO(un9_6_0_cry_38));
  XORCY un9_6_0_s_37(.LI(un9_6_0_axb_37),.CI(un9_6_0_cry_36),.O(un9_6[37:37]));
  MUXCY_L un9_6_0_cry_37_cZ(.DI(un9_11[37:37]),.CI(un9_6_0_cry_36),.S(un9_6_0_axb_37),.LO(un9_6_0_cry_37));
  XORCY un9_6_0_s_36(.LI(un9_6_0_axb_36),.CI(un9_6_0_cry_35),.O(un9_6[36:36]));
  MUXCY_L un9_6_0_cry_36_cZ(.DI(un9_6_0_cry_36_RNO),.CI(un9_6_0_cry_35),.S(un9_6_0_axb_36),.LO(un9_6_0_cry_36));
  XORCY un9_6_0_s_35(.LI(un9_6_0_axb_35),.CI(un9_6_0_cry_34),.O(un9_6[35:35]));
  MUXCY_L un9_6_0_cry_35_cZ(.DI(un9_6_0_cry_35_RNO),.CI(un9_6_0_cry_34),.S(un9_6_0_axb_35),.LO(un9_6_0_cry_35));
  XORCY un9_6_0_s_34(.LI(un9_6_0_axb_34),.CI(un9_6_0_cry_33),.O(un9_6[34:34]));
  MUXCY_L un9_6_0_cry_34_cZ(.DI(un9_6_0_cry_34_RNO),.CI(un9_6_0_cry_33),.S(un9_6_0_axb_34),.LO(un9_6_0_cry_34));
  XORCY un9_6_0_s_33(.LI(un9_6_0_axb_33),.CI(un9_6_0_cry_32),.O(un9_6[33:33]));
  MUXCY_L un9_6_0_cry_33_cZ(.DI(un9_6_0_cry_33_RNO),.CI(un9_6_0_cry_32),.S(un9_6_0_axb_33),.LO(un9_6_0_cry_33));
  XORCY un9_6_0_s_32(.LI(un9_6_0_axb_32),.CI(un9_6_0_cry_31),.O(un9_6[32:32]));
  MUXCY_L un9_6_0_cry_32_cZ(.DI(un9_6_0_cry_32_RNO),.CI(un9_6_0_cry_31),.S(un9_6_0_axb_32),.LO(un9_6_0_cry_32));
  XORCY un9_6_0_s_31(.LI(un9_6_0_axb_31),.CI(un9_6_0_cry_30),.O(un9_6[31:31]));
  MUXCY_L un9_6_0_cry_31_cZ(.DI(un9_6_0_cry_31_RNO),.CI(un9_6_0_cry_30),.S(un9_6_0_axb_31),.LO(un9_6_0_cry_31));
  XORCY un9_6_0_s_30(.LI(un9_6_0_axb_30),.CI(un9_6_0_cry_29),.O(un9_6[30:30]));
  MUXCY_L un9_6_0_cry_30_cZ(.DI(un9_6_0_cry_30_RNO),.CI(un9_6_0_cry_29),.S(un9_6_0_axb_30),.LO(un9_6_0_cry_30));
  XORCY un9_6_0_s_29(.LI(un9_6_0_axb_29),.CI(un9_6_0_cry_28),.O(un9_6[29:29]));
  MUXCY_L un9_6_0_cry_29_cZ(.DI(un9_6_0_cry_29_RNO),.CI(un9_6_0_cry_28),.S(un9_6_0_axb_29),.LO(un9_6_0_cry_29));
  XORCY un9_6_0_s_28(.LI(un9_6_0_axb_28),.CI(un9_6_0_cry_27),.O(un9_6[28:28]));
  MUXCY_L un9_6_0_cry_28_cZ(.DI(un9_6_0_cry_28_RNO),.CI(un9_6_0_cry_27),.S(un9_6_0_axb_28),.LO(un9_6_0_cry_28));
  XORCY un9_6_0_s_27(.LI(un9_6_0_axb_27),.CI(un9_6_0_cry_26),.O(un9_6[27:27]));
  MUXCY_L un9_6_0_cry_27_cZ(.DI(un9_6_0_cry_27_RNO),.CI(un9_6_0_cry_26),.S(un9_6_0_axb_27),.LO(un9_6_0_cry_27));
  XORCY un9_6_0_s_26(.LI(un9_6_0_axb_26),.CI(un9_6_0_cry_25),.O(un9_6[26:26]));
  MUXCY_L un9_6_0_cry_26_cZ(.DI(un9_6_0_cry_26_RNO),.CI(un9_6_0_cry_25),.S(un9_6_0_axb_26),.LO(un9_6_0_cry_26));
  XORCY un9_6_0_s_25(.LI(un9_6_0_axb_25),.CI(un9_6_0_cry_24),.O(un9_6[25:25]));
  MUXCY_L un9_6_0_cry_25_cZ(.DI(un9_6_0_cry_25_RNO),.CI(un9_6_0_cry_24),.S(un9_6_0_axb_25),.LO(un9_6_0_cry_25));
  XORCY un9_6_0_s_24(.LI(un9_6_0_axb_24),.CI(un9_6_0_cry_23),.O(un9_6[24:24]));
  MUXCY_L un9_6_0_cry_24_cZ(.DI(un9_6_0_cry_24_RNO),.CI(un9_6_0_cry_23),.S(un9_6_0_axb_24),.LO(un9_6_0_cry_24));
  XORCY un9_6_0_s_23(.LI(un9_6_0_axb_23),.CI(un9_6_0_cry_22),.O(un9_6[23:23]));
  MUXCY_L un9_6_0_cry_23_cZ(.DI(un9_6_0_cry_23_RNO),.CI(un9_6_0_cry_22),.S(un9_6_0_axb_23),.LO(un9_6_0_cry_23));
  XORCY un9_6_0_s_22(.LI(un9_6_0_axb_22),.CI(un9_6_0_cry_21),.O(un9_6[22:22]));
  MUXCY_L un9_6_0_cry_22_cZ(.DI(un9_6_0_cry_22_RNO),.CI(un9_6_0_cry_21),.S(un9_6_0_axb_22),.LO(un9_6_0_cry_22));
  XORCY un9_6_0_s_21(.LI(un9_6_0_axb_21),.CI(un9_6_0_cry_20),.O(un9_6[21:21]));
  MUXCY_L un9_6_0_cry_21_cZ(.DI(ZFF_Y1_9_rep1),.CI(un9_6_0_cry_20),.S(un9_6_0_axb_21),.LO(un9_6_0_cry_21));
  XORCY un9_6_0_s_20(.LI(un9_6_0_axb_20),.CI(un9_6_0_cry_19),.O(un9_6[20:20]));
  MUXCY_L un9_6_0_cry_20_cZ(.DI(un9_6_0_cry_20_RNO),.CI(un9_6_0_cry_19),.S(un9_6_0_axb_20),.LO(un9_6_0_cry_20));
  XORCY un9_6_0_s_19(.LI(un9_6_0_axb_19),.CI(un9_6_0_cry_18),.O(un9_6[19:19]));
  MUXCY_L un9_6_0_cry_19_cZ(.DI(un9_6_0_cry_19_RNO),.CI(un9_6_0_cry_18),.S(un9_6_0_axb_19),.LO(un9_6_0_cry_19));
  XORCY un9_6_0_s_18(.LI(un9_6_0_axb_18),.CI(un9_6_0_cry_17),.O(un9_6[18:18]));
  MUXCY_L un9_6_0_cry_18_cZ(.DI(un9_6_0_cry_18_RNO),.CI(un9_6_0_cry_17),.S(un9_6_0_axb_18),.LO(un9_6_0_cry_18));
  XORCY un9_6_0_s_17(.LI(un9_6_0_axb_17),.CI(un9_6_0_cry_16),.O(un9_6[17:17]));
  MUXCY_L un9_6_0_cry_17_cZ(.DI(un9_6_0_cry_17_RNO),.CI(un9_6_0_cry_16),.S(un9_6_0_axb_17),.LO(un9_6_0_cry_17));
  XORCY un9_6_0_s_16(.LI(un9_6_0_axb_16),.CI(un9_6_0_cry_15),.O(un9_6[16:16]));
  MUXCY_L un9_6_0_cry_16_cZ(.DI(un9_6_0_cry_16_RNO),.CI(un9_6_0_cry_15),.S(un9_6_0_axb_16),.LO(un9_6_0_cry_16));
  XORCY un9_6_0_s_15(.LI(un9_6_0_axb_15),.CI(un9_6_0_cry_14),.O(un9_6[15:15]));
  MUXCY_L un9_6_0_cry_15_cZ(.DI(un9_6_0_cry_15_RNO),.CI(un9_6_0_cry_14),.S(un9_6_0_axb_15),.LO(un9_6_0_cry_15));
  XORCY un9_6_0_s_14(.LI(un9_6_0_axb_14),.CI(un9_6_0_cry_13),.O(un9_6[14:14]));
  MUXCY_L un9_6_0_cry_14_cZ(.DI(un9_6_0_cry_14_RNO),.CI(un9_6_0_cry_13),.S(un9_6_0_axb_14),.LO(un9_6_0_cry_14));
  XORCY un9_6_0_s_13(.LI(un9_6_0_axb_13),.CI(un9_6_0_cry_12),.O(un9_6[13:13]));
  MUXCY_L un9_6_0_cry_13_cZ(.DI(un9_6_0_cry_13_RNO),.CI(un9_6_0_cry_12),.S(un9_6_0_axb_13),.LO(un9_6_0_cry_13));
  XORCY un9_6_0_s_12(.LI(un9_6_0_axb_12),.CI(un9_6_0_cry_11),.O(un9_6[12:12]));
  MUXCY_L un9_6_0_cry_12_cZ(.DI(un9_6_0_cry_12_RNO),.CI(un9_6_0_cry_11),.S(un9_6_0_axb_12),.LO(un9_6_0_cry_12));
  XORCY un9_6_0_s_11(.LI(un9_6_0_axb_11),.CI(un9_6_0_cry_10),.O(un9_6[11:11]));
  MUXCY_L un9_6_0_cry_11_cZ(.DI(un9_6_0_cry_11_RNO),.CI(un9_6_0_cry_10),.S(un9_6_0_axb_11),.LO(un9_6_0_cry_11));
  XORCY un9_6_0_s_10(.LI(un9_6_0_axb_10),.CI(un9_6_0_cry_9),.O(un9_6[10:10]));
  MUXCY_L un9_6_0_cry_10_cZ(.DI(GND),.CI(un9_6_0_cry_9),.S(un9_6_0_axb_10),.LO(un9_6_0_cry_10));
  MUXCY_L un9_6_0_cry_9_cZ(.DI(GND),.CI(un9_6_0_cry_8),.S(un9_6_0_cry_9_RNO),.LO(un9_6_0_cry_9));
  XORCY un9_6_0_s_8(.LI(un9_6_0_axb_8),.CI(un9_6_0_cry_7),.O(un9_6[8:8]));
  XORCY un9_6_0_s_7(.LI(un9_6_0_axb_7),.CI(un9_6_0_cry_6),.O(un9_6[7:7]));
  MUXCY_L un9_6_0_cry_7_cZ(.DI(un9_6_0_cry_7_RNO),.CI(un9_6_0_cry_6),.S(un9_6_0_axb_7),.LO(un9_6_0_cry_7));
  XORCY un9_6_0_s_6(.LI(un9_6_0_axb_6),.CI(un9_6_0_cry_5),.O(un9_6[6:6]));
  MUXCY_L un9_6_0_cry_6_cZ(.DI(un9_6_0_cry_6_RNO),.CI(un9_6_0_cry_5),.S(un9_6_0_axb_6),.LO(un9_6_0_cry_6));
  MUXCY_L un9_6_0_cry_5_cZ(.DI(un9_6_0_cry_5_RNO),.CI(GND),.S(un9_6_0_cry_5_RNO_0),.LO(un9_6_0_cry_5));
  XORCY un9_s_45_cZ(.LI(un9_axb_45),.CI(un9_cry_44),.O(un9_s_45));
  XORCY un9_s_44_cZ(.LI(un9_axb_44),.CI(un9_cry_43),.O(un9_s_44));
  MUXCY_L un9_cry_44_cZ(.DI(un9_cry_44_RNO),.CI(un9_cry_43),.S(un9_axb_44),.LO(un9_cry_44));
  XORCY un9_s_43_cZ(.LI(un9_axb_43),.CI(un9_cry_42),.O(un9_s_43));
  MUXCY_L un9_cry_43_cZ(.DI(un9_cry_43_RNO),.CI(un9_cry_42),.S(un9_axb_43),.LO(un9_cry_43));
  XORCY un9_s_42_cZ(.LI(un9_axb_42),.CI(un9_cry_41),.O(un9_s_42));
  MUXCY_L un9_cry_42_cZ(.DI(un9_cry_42_RNO),.CI(un9_cry_41),.S(un9_axb_42),.LO(un9_cry_42));
  XORCY un9_s_41_cZ(.LI(un9_axb_41),.CI(un9_cry_40),.O(un9_s_41));
  MUXCY_L un9_cry_41_cZ(.DI(un9_cry_41_RNO),.CI(un9_cry_40),.S(un9_axb_41),.LO(un9_cry_41));
  XORCY un9_s_40_cZ(.LI(un9_axb_40),.CI(un9_cry_39),.O(un9_s_40));
  MUXCY_L un9_cry_40_cZ(.DI(un9_o5_39),.CI(un9_cry_39),.S(un9_axb_40),.LO(un9_cry_40));
  XORCY un9_s_39_cZ(.LI(un9_axb_39),.CI(un9_cry_38),.O(un9_s_39));
  MUXCY_L un9_cry_39_cZ(.DI(un9_o5_38),.CI(un9_cry_38),.S(un9_axb_39),.LO(un9_cry_39));
  XORCY un9_s_38_cZ(.LI(un9_axb_38),.CI(un9_cry_37),.O(un9_s_38));
  MUXCY_L un9_cry_38_cZ(.DI(un9_o5_37),.CI(un9_cry_37),.S(un9_axb_38),.LO(un9_cry_38));
  XORCY un9_s_37_cZ(.LI(un9_axb_37),.CI(un9_cry_36),.O(un9_s_37));
  MUXCY_L un9_cry_37_cZ(.DI(un9_o5_36),.CI(un9_cry_36),.S(un9_axb_37),.LO(un9_cry_37));
  XORCY un9_s_36_cZ(.LI(un9_axb_36),.CI(un9_cry_35),.O(un9_s_36));
  MUXCY_L un9_cry_36_cZ(.DI(un9_o5_35),.CI(un9_cry_35),.S(un9_axb_36),.LO(un9_cry_36));
  XORCY un9_s_35_cZ(.LI(un9_axb_35),.CI(un9_cry_34),.O(un9_s_35));
  MUXCY_L un9_cry_35_cZ(.DI(un9_o5_34),.CI(un9_cry_34),.S(un9_axb_35),.LO(un9_cry_35));
  XORCY un9_s_34_cZ(.LI(un9_axb_34),.CI(un9_cry_33),.O(un9_s_34));
  MUXCY_L un9_cry_34_cZ(.DI(un9_o5_33),.CI(un9_cry_33),.S(un9_axb_34),.LO(un9_cry_34));
  XORCY un9_s_33_cZ(.LI(un9_axb_33),.CI(un9_cry_32),.O(un9_s_33));
  MUXCY_L un9_cry_33_cZ(.DI(un9_o5_32),.CI(un9_cry_32),.S(un9_axb_33),.LO(un9_cry_33));
  XORCY un9_s_32_cZ(.LI(un9_axb_32),.CI(un9_cry_31),.O(un9_s_32));
  MUXCY_L un9_cry_32_cZ(.DI(un9_o5_31),.CI(un9_cry_31),.S(un9_axb_32),.LO(un9_cry_32));
  XORCY un9_s_31_cZ(.LI(un9_axb_31),.CI(un9_cry_30),.O(un9_s_31));
  MUXCY_L un9_cry_31_cZ(.DI(un9_o5_30),.CI(un9_cry_30),.S(un9_axb_31),.LO(un9_cry_31));
  XORCY un9_s_30_cZ(.LI(un9_axb_30),.CI(un9_cry_29),.O(un9_s_30));
  MUXCY_L un9_cry_30_cZ(.DI(un9_o5_29),.CI(un9_cry_29),.S(un9_axb_30),.LO(un9_cry_30));
  XORCY un9_s_29_cZ(.LI(un9_axb_29),.CI(un9_cry_28),.O(un9_s_29));
  MUXCY_L un9_cry_29_cZ(.DI(un9_o5_28),.CI(un9_cry_28),.S(un9_axb_29),.LO(un9_cry_29));
  XORCY un9_s_28_cZ(.LI(un9_axb_28),.CI(un9_cry_27),.O(un9_s_28));
  MUXCY_L un9_cry_28_cZ(.DI(un9_o5_27),.CI(un9_cry_27),.S(un9_axb_28),.LO(un9_cry_28));
  MUXCY_L un9_cry_27_cZ(.DI(un9_o5_26),.CI(un9_cry_26),.S(un9_axb_27),.LO(un9_cry_27));
  MUXCY_L un9_cry_26_cZ(.DI(un9_o5_25),.CI(un9_cry_25),.S(un9_axb_26),.LO(un9_cry_26));
  MUXCY_L un9_cry_25_cZ(.DI(un9_o5_24),.CI(un9_cry_24),.S(un9_axb_25),.LO(un9_cry_25));
  MUXCY_L un9_cry_24_cZ(.DI(un9_o5_23),.CI(un9_cry_23),.S(un9_axb_24),.LO(un9_cry_24));
  MUXCY_L un9_cry_23_cZ(.DI(un9_o5_22),.CI(un9_cry_22),.S(un9_axb_23),.LO(un9_cry_23));
  MUXCY_L un9_cry_22_cZ(.DI(un9_o5_21),.CI(un9_cry_21),.S(un9_axb_22),.LO(un9_cry_22));
  MUXCY_L un9_cry_21_cZ(.DI(un9_o5_20),.CI(un9_cry_20),.S(un9_axb_21),.LO(un9_cry_21));
  MUXCY_L un9_cry_20_cZ(.DI(un9_o5_19),.CI(un9_cry_19),.S(un9_axb_20),.LO(un9_cry_20));
  MUXCY_L un9_cry_19_cZ(.DI(un9_o5_18),.CI(un9_cry_18),.S(un9_axb_19),.LO(un9_cry_19));
  MUXCY_L un9_cry_18_cZ(.DI(un9_o5_17),.CI(un9_cry_17),.S(un9_axb_18),.LO(un9_cry_18));
  MUXCY_L un9_cry_17_cZ(.DI(un9_o5_16),.CI(un9_cry_16),.S(un9_axb_17),.LO(un9_cry_17));
  MUXCY_L un9_cry_16_cZ(.DI(un9_o5_15),.CI(un9_cry_15),.S(un9_axb_16),.LO(un9_cry_16));
  MUXCY_L un9_cry_15_cZ(.DI(un9_o5_14),.CI(un9_cry_14),.S(un9_axb_15),.LO(un9_cry_15));
  MUXCY_L un9_cry_14_cZ(.DI(un9_o5_13),.CI(un9_cry_13),.S(un9_axb_14),.LO(un9_cry_14));
  MUXCY_L un9_cry_13_cZ(.DI(un9_o5_12),.CI(un9_cry_12),.S(un9_axb_13),.LO(un9_cry_13));
  MUXCY_L un9_cry_12_cZ(.DI(un9_o5_11),.CI(un9_cry_11),.S(un9_axb_12),.LO(un9_cry_12));
  MUXCY_L un9_cry_11_cZ(.DI(un9_o5_10),.CI(un9_cry_10),.S(un9_axb_11),.LO(un9_cry_11));
  MUXCY_L un9_cry_10_cZ(.DI(un9_o5_9),.CI(un9_cry_9),.S(un9_axb_10),.LO(un9_cry_10));
  MUXCY_L un9_cry_9_cZ(.DI(un9_o5_8),.CI(un9_cry_8),.S(un9_axb_9),.LO(un9_cry_9));
  MUXCY_L un9_cry_8_cZ(.DI(un9_o5_7),.CI(un9_cry_7),.S(un9_axb_8),.LO(un9_cry_8));
  MUXCY_L un9_cry_7_cZ(.DI(un9_cry_7_RNO),.CI(un9_cry_6),.S(un9_axb_7),.LO(un9_cry_7));
  MUXCY_L un9_cry_6_cZ(.DI(un9_6[8:8]),.CI(un9_cry_5),.S(un9_axb_6),.LO(un9_cry_6));
  MUXCY_L un9_cry_5_cZ(.DI(un9_6[7:7]),.CI(un9_cry_4),.S(un9_axb_5),.LO(un9_cry_5));
  MUXCY_L un9_cry_4_cZ(.DI(un9_6[6:6]),.CI(un9_cry_3),.S(un9_axb_4),.LO(un9_cry_4));
  MUXCY_L un9_cry_3_cZ(.DI(un9_6[5:5]),.CI(un9_cry_2),.S(un9_axb_3),.LO(un9_cry_3));
  MUXCY_L un9_cry_2_cZ(.DI(un9_6[4:4]),.CI(un9_cry_1),.S(un9_axb_2),.LO(un9_cry_2));
  MUXCY_L un9_cry_1_cZ(.DI(un9_6[3:3]),.CI(un9_cry_0),.S(un9_axb_1),.LO(un9_cry_1));
  MUXCY_L un9_cry_0_cZ(.DI(VCC),.CI(un9_cry_0_cy),.S(un9_6[2:2]),.LO(un9_cry_0));
  XORCY Y_out_double_2_6_0_s_17(.LI(Y_out_double_2_6_0_axb_17),.CI(Y_out_double_2_6_0_cry_16),.O(Y_out_double_2_6[17:17]));
  XORCY Y_out_double_2_6_0_s_16(.LI(Y_out_double_2_6_0_axb_16),.CI(Y_out_double_2_6_0_cry_15),.O(Y_out_double_2_6[16:16]));
  MUXCY_L Y_out_double_2_6_0_cry_16_cZ(.DI(Y_out_double_2_6_0_o5_15),.CI(Y_out_double_2_6_0_cry_15),.S(Y_out_double_2_6_0_axb_16),.LO(Y_out_double_2_6_0_cry_16));
  XORCY Y_out_double_2_6_0_s_15(.LI(Y_out_double_2_6_0_axb_15),.CI(Y_out_double_2_6_0_cry_14),.O(Y_out_double_2_6[15:15]));
  MUXCY_L Y_out_double_2_6_0_cry_15_cZ(.DI(Y_out_double_2_6_0_o5_14),.CI(Y_out_double_2_6_0_cry_14),.S(Y_out_double_2_6_0_axb_15),.LO(Y_out_double_2_6_0_cry_15));
  XORCY Y_out_double_2_6_0_s_14(.LI(Y_out_double_2_6_0_axb_14),.CI(Y_out_double_2_6_0_cry_13),.O(Y_out_double_2_6[14:14]));
  MUXCY_L Y_out_double_2_6_0_cry_14_cZ(.DI(Y_out_double_2_6_0_o5_13),.CI(Y_out_double_2_6_0_cry_13),.S(Y_out_double_2_6_0_axb_14),.LO(Y_out_double_2_6_0_cry_14));
  XORCY Y_out_double_2_6_0_s_13(.LI(Y_out_double_2_6_0_axb_13),.CI(Y_out_double_2_6_0_cry_12),.O(Y_out_double_2_6[13:13]));
  MUXCY_L Y_out_double_2_6_0_cry_13_cZ(.DI(Y_out_double_2_6_0_o5_12),.CI(Y_out_double_2_6_0_cry_12),.S(Y_out_double_2_6_0_axb_13),.LO(Y_out_double_2_6_0_cry_13));
  XORCY Y_out_double_2_6_0_s_12(.LI(Y_out_double_2_6_0_axb_12),.CI(Y_out_double_2_6_0_cry_11),.O(Y_out_double_2_6[12:12]));
  MUXCY_L Y_out_double_2_6_0_cry_12_cZ(.DI(Y_out_double_2_6_0_o5_11),.CI(Y_out_double_2_6_0_cry_11),.S(Y_out_double_2_6_0_axb_12),.LO(Y_out_double_2_6_0_cry_12));
  XORCY Y_out_double_2_6_0_s_11(.LI(Y_out_double_2_6_0_axb_11),.CI(Y_out_double_2_6_0_cry_10),.O(Y_out_double_2_6[11:11]));
  MUXCY_L Y_out_double_2_6_0_cry_11_cZ(.DI(Y_out_double_2_6_0_o5_10),.CI(Y_out_double_2_6_0_cry_10),.S(Y_out_double_2_6_0_axb_11),.LO(Y_out_double_2_6_0_cry_11));
  XORCY Y_out_double_2_6_0_s_10(.LI(Y_out_double_2_6_0_axb_10),.CI(Y_out_double_2_6_0_cry_9),.O(Y_out_double_2_6[10:10]));
  MUXCY_L Y_out_double_2_6_0_cry_10_cZ(.DI(Y_out_double_2_6_0_o5_9),.CI(Y_out_double_2_6_0_cry_9),.S(Y_out_double_2_6_0_axb_10),.LO(Y_out_double_2_6_0_cry_10));
  XORCY Y_out_double_2_6_0_s_9(.LI(Y_out_double_2_6_0_axb_9),.CI(Y_out_double_2_6_0_cry_8),.O(Y_out_double_2_6[9:9]));
  MUXCY_L Y_out_double_2_6_0_cry_9_cZ(.DI(Y_out_double_2_6_0_o5_8),.CI(Y_out_double_2_6_0_cry_8),.S(Y_out_double_2_6_0_axb_9),.LO(Y_out_double_2_6_0_cry_9));
  XORCY Y_out_double_2_6_0_s_8(.LI(Y_out_double_2_6_0_axb_8),.CI(Y_out_double_2_6_0_cry_7),.O(Y_out_double_2_6[8:8]));
  MUXCY_L Y_out_double_2_6_0_cry_8_cZ(.DI(Y_out_double_2_6_0_o5_7),.CI(Y_out_double_2_6_0_cry_7),.S(Y_out_double_2_6_0_axb_8),.LO(Y_out_double_2_6_0_cry_8));
  XORCY Y_out_double_2_6_0_s_7(.LI(Y_out_double_2_6_0_axb_7),.CI(Y_out_double_2_6_0_cry_6),.O(Y_out_double_2_6[7:7]));
  MUXCY_L Y_out_double_2_6_0_cry_7_cZ(.DI(Y_out_double_2_6_0_o5_6),.CI(Y_out_double_2_6_0_cry_6),.S(Y_out_double_2_6_0_axb_7),.LO(Y_out_double_2_6_0_cry_7));
  XORCY Y_out_double_2_6_0_s_6(.LI(Y_out_double_2_6_0_axb_6),.CI(Y_out_double_2_6_0_cry_5),.O(Y_out_double_2_6[6:6]));
  MUXCY_L Y_out_double_2_6_0_cry_6_cZ(.DI(Y_out_double_2_6_0_o5_5),.CI(Y_out_double_2_6_0_cry_5),.S(Y_out_double_2_6_0_axb_6),.LO(Y_out_double_2_6_0_cry_6));
  XORCY Y_out_double_2_6_0_s_5(.LI(Y_out_double_2_6_0_axb_5),.CI(Y_out_double_2_6_0_cry_4),.O(Y_out_double_2_6[5:5]));
  MUXCY_L Y_out_double_2_6_0_cry_5_cZ(.DI(Y_out_double_2_6_0_o5_4),.CI(Y_out_double_2_6_0_cry_4),.S(Y_out_double_2_6_0_axb_5),.LO(Y_out_double_2_6_0_cry_5));
  XORCY Y_out_double_2_6_0_s_4(.LI(Y_out_double_2_6_0_axb_4),.CI(Y_out_double_2_6_0_cry_3),.O(Y_out_double_2_6[4:4]));
  MUXCY_L Y_out_double_2_6_0_cry_4_cZ(.DI(Y_out_double_2_6_0_o5_3),.CI(Y_out_double_2_6_0_cry_3),.S(Y_out_double_2_6_0_axb_4),.LO(Y_out_double_2_6_0_cry_4));
  XORCY Y_out_double_2_6_0_s_3(.LI(Y_out_double_2_6_0_axb_3),.CI(Y_out_double_2_6_0_cry_2),.O(Y_out_double_2_6[3:3]));
  MUXCY_L Y_out_double_2_6_0_cry_3_cZ(.DI(Y_out_double_2_6_0_o5_2),.CI(Y_out_double_2_6_0_cry_2),.S(Y_out_double_2_6_0_axb_3),.LO(Y_out_double_2_6_0_cry_3));
  XORCY Y_out_double_2_6_0_s_2(.LI(Y_out_double_2_6_0_axb_2),.CI(Y_out_double_2_6_0_cry_1),.O(Y_out_double_2_6[2:2]));
  MUXCY_L Y_out_double_2_6_0_cry_2_cZ(.DI(Y_out_double_2_6_0_o5_1),.CI(Y_out_double_2_6_0_cry_1),.S(Y_out_double_2_6_0_axb_2),.LO(Y_out_double_2_6_0_cry_2));
  XORCY Y_out_double_2_6_0_s_1(.LI(Y_out_double_2_6_0_axb_1),.CI(Y_out_double_2_6_0_cry_0),.O(Y_out_double_2_6[1:1]));
  MUXCY_L Y_out_double_2_6_0_cry_1_cZ(.DI(GND),.CI(Y_out_double_2_6_0_cry_0),.S(Y_out_double_2_6_0_axb_1),.LO(Y_out_double_2_6_0_cry_1));
  XORCY Y_out_double_2_6_0_s_0(.LI(Y_out_double_2_6_0_axb_0),.CI(pgZFF_X1[0:0]),.O(Y_out_double_2_6[0:0]));
  MUXCY_L Y_out_double_2_6_0_cry_0_cZ(.DI(pgZFF_Y1_i),.CI(pgZFF_X1[0:0]),.S(Y_out_double_2_6_0_axb_0),.LO(Y_out_double_2_6_0_cry_0));
  XORCY un6_0_6_s_22(.LI(un6_0_6_axb_22),.CI(un6_0_6_cry_21),.O(un6_0_6[27:27]));
  MUXCY un6_0_6_cry_22(.DI(GND),.CI(un6_0_6_cry_21),.S(un6_0_6_axb_22),.O(un6_0_6_0[28:28]));
  XORCY un6_0_6_s_21(.LI(un6_0_6_axb_21),.CI(un6_0_6_cry_20),.O(un6_0_6[26:26]));
  MUXCY_L un6_0_6_cry_21_cZ(.DI(un6_0_6_43),.CI(un6_0_6_cry_20),.S(un6_0_6_axb_21),.LO(un6_0_6_cry_21));
  XORCY un6_0_6_s_20(.LI(un6_0_6_axb_20),.CI(un6_0_6_cry_19),.O(un6_0_6[25:25]));
  MUXCY_L un6_0_6_cry_20_cZ(.DI(un6_0_6_cry_20_RNO),.CI(un6_0_6_cry_19),.S(un6_0_6_axb_20),.LO(un6_0_6_cry_20));
  XORCY un6_0_6_s_19(.LI(un6_0_6_axb_19),.CI(un6_0_6_cry_18),.O(un6_0_6[24:24]));
  MUXCY_L un6_0_6_cry_19_cZ(.DI(un6_0_6_cry_19_RNO),.CI(un6_0_6_cry_18),.S(un6_0_6_axb_19),.LO(un6_0_6_cry_19));
  XORCY un6_0_6_s_18(.LI(un6_0_6_axb_18),.CI(un6_0_6_cry_17),.O(un6_0_6[23:23]));
  MUXCY_L un6_0_6_cry_18_cZ(.DI(un6_0_6_cry_18_RNO),.CI(un6_0_6_cry_17),.S(un6_0_6_axb_18),.LO(un6_0_6_cry_18));
  XORCY un6_0_6_s_17(.LI(un6_0_6_axb_17),.CI(un6_0_6_cry_16),.O(un6_0_6[22:22]));
  MUXCY_L un6_0_6_cry_17_cZ(.DI(un6_0_6_cry_17_RNO),.CI(un6_0_6_cry_16),.S(un6_0_6_axb_17),.LO(un6_0_6_cry_17));
  XORCY un6_0_6_s_16(.LI(un6_0_6_axb_16),.CI(un6_0_6_cry_15),.O(un6_0_6[21:21]));
  MUXCY_L un6_0_6_cry_16_cZ(.DI(un6_0_6_cry_16_RNO),.CI(un6_0_6_cry_15),.S(un6_0_6_axb_16),.LO(un6_0_6_cry_16));
  XORCY un6_0_6_s_15(.LI(un6_0_6_axb_15),.CI(un6_0_6_cry_14),.O(un6_0_6[20:20]));
  MUXCY_L un6_0_6_cry_15_cZ(.DI(un6_0_6_cry_15_RNO),.CI(un6_0_6_cry_14),.S(un6_0_6_axb_15),.LO(un6_0_6_cry_15));
  XORCY un6_0_6_s_14(.LI(un6_0_6_axb_14),.CI(un6_0_6_cry_13),.O(un6_0_6[19:19]));
  MUXCY_L un6_0_6_cry_14_cZ(.DI(un6_0_6_cry_14_RNO),.CI(un6_0_6_cry_13),.S(un6_0_6_axb_14),.LO(un6_0_6_cry_14));
  XORCY un6_0_6_s_13(.LI(un6_0_6_axb_13),.CI(un6_0_6_cry_12),.O(un6_0_6[18:18]));
  MUXCY_L un6_0_6_cry_13_cZ(.DI(un6_0_6_cry_13_RNO),.CI(un6_0_6_cry_12),.S(un6_0_6_axb_13),.LO(un6_0_6_cry_13));
  XORCY un6_0_6_s_12(.LI(un6_0_6_axb_12),.CI(un6_0_6_cry_11),.O(un6_0_6[17:17]));
  MUXCY_L un6_0_6_cry_12_cZ(.DI(un6_0_6_cry_12_RNO),.CI(un6_0_6_cry_11),.S(un6_0_6_axb_12),.LO(un6_0_6_cry_12));
  XORCY un6_0_6_s_11(.LI(un6_0_6_axb_11),.CI(un6_0_6_cry_10),.O(un6_0_6[16:16]));
  MUXCY_L un6_0_6_cry_11_cZ(.DI(un6_0_6_cry_11_RNO),.CI(un6_0_6_cry_10),.S(un6_0_6_axb_11),.LO(un6_0_6_cry_11));
  XORCY un6_0_6_s_10(.LI(un6_0_6_axb_10),.CI(un6_0_6_cry_9),.O(un6_0_6[15:15]));
  MUXCY_L un6_0_6_cry_10_cZ(.DI(un6_0_6_cry_10_RNO),.CI(un6_0_6_cry_9),.S(un6_0_6_axb_10),.LO(un6_0_6_cry_10));
  XORCY un6_0_6_s_9(.LI(un6_0_6_axb_9),.CI(un6_0_6_cry_8),.O(un6_0_6[14:14]));
  MUXCY_L un6_0_6_cry_9_cZ(.DI(un6_0_6_cry_9_RNO),.CI(un6_0_6_cry_8),.S(un6_0_6_axb_9),.LO(un6_0_6_cry_9));
  XORCY un6_0_6_s_8(.LI(un6_0_6_axb_8),.CI(un6_0_6_cry_7),.O(un6_0_6[13:13]));
  MUXCY_L un6_0_6_cry_8_cZ(.DI(un6_0_6_cry_8_RNO),.CI(un6_0_6_cry_7),.S(un6_0_6_axb_8),.LO(un6_0_6_cry_8));
  XORCY un6_0_6_s_7(.LI(un6_0_6_axb_7),.CI(un6_0_6_cry_6),.O(un6_0_6[12:12]));
  MUXCY_L un6_0_6_cry_7_cZ(.DI(un6_0_6_cry_7_RNO),.CI(un6_0_6_cry_6),.S(un6_0_6_axb_7),.LO(un6_0_6_cry_7));
  XORCY un6_0_6_s_6(.LI(un6_0_6_axb_6),.CI(un6_0_6_cry_5),.O(un6_0_6[11:11]));
  MUXCY_L un6_0_6_cry_6_cZ(.DI(un6_0_6_cry_6_RNO),.CI(un6_0_6_cry_5),.S(un6_0_6_axb_6),.LO(un6_0_6_cry_6));
  XORCY un6_0_6_s_5(.LI(un6_0_6_axb_5),.CI(un6_0_6_cry_4),.O(un6_0_6[10:10]));
  MUXCY_L un6_0_6_cry_5_cZ(.DI(un6_0_6_cry_5_RNO),.CI(un6_0_6_cry_4),.S(un6_0_6_axb_5),.LO(un6_0_6_cry_5));
  XORCY un6_0_6_s_4(.LI(un6_0_6_axb_4),.CI(un6_0_6_cry_3),.O(un6_0_6[9:9]));
  MUXCY_L un6_0_6_cry_4_cZ(.DI(un6_0_6_cry_4_RNO),.CI(un6_0_6_cry_3),.S(un6_0_6_axb_4),.LO(un6_0_6_cry_4));
  XORCY un6_0_6_s_3(.LI(un6_0_6_axb_3),.CI(un6_0_6_cry_2),.O(un6_0_6[8:8]));
  MUXCY_L un6_0_6_cry_3_cZ(.DI(N_2372_i),.CI(un6_0_6_cry_2),.S(un6_0_6_axb_3),.LO(un6_0_6_cry_3));
  XORCY un6_0_6_s_2(.LI(un6_0_6_axb_2),.CI(un6_0_6_cry_1),.O(un6_0_6[7:7]));
  MUXCY_L un6_0_6_cry_2_cZ(.DI(ZFF_X0[0:0]),.CI(un6_0_6_cry_1),.S(un6_0_6_axb_2),.LO(un6_0_6_cry_2));
  XORCY un6_0_6_s_1(.LI(un6_0_6_axb_1),.CI(un6_0_6_cry_0),.O(un6_0_6[6:6]));
  MUXCY_L un6_0_6_cry_1_cZ(.DI(ZFF_X0_1_rep1),.CI(un6_0_6_cry_0),.S(un6_0_6_axb_1),.LO(un6_0_6_cry_1));
  MUXCY_L un6_0_6_cry_0_cZ(.DI(N_2379_i),.CI(GND),.S(un6_0_6_cry_0_sf),.LO(un6_0_6_cry_0));
  XORCY un6_0_0_s_43_cZ(.LI(un6_0_0_axb_43),.CI(un6_0_0_cry_42),.O(un6_0_0_s_43));
  XORCY un6_0_0_s_42_cZ(.LI(un6_0_0_axb_42),.CI(un6_0_0_cry_41),.O(un6_0_0_s_42));
  MUXCY_L un6_0_0_cry_42_cZ(.DI(un6_0_0_o5_41),.CI(un6_0_0_cry_41),.S(un6_0_0_axb_42),.LO(un6_0_0_cry_42));
  XORCY un6_0_0_s_41_cZ(.LI(un6_0_0_axb_41),.CI(un6_0_0_cry_40),.O(un6_0_0_s_41));
  MUXCY_L un6_0_0_cry_41_cZ(.DI(GND),.CI(un6_0_0_cry_40),.S(un6_0_0_axb_41),.LO(un6_0_0_cry_41));
  XORCY un6_0_0_s_40_cZ(.LI(N_2007_i),.CI(un6_0_0_cry_39),.O(un6_0_0_s_40));
  MUXCY_L un6_0_0_cry_40_cZ(.DI(VCC),.CI(un6_0_0_cry_39),.S(N_2007_i),.LO(un6_0_0_cry_40));
  XORCY un6_0_0_s_39_cZ(.LI(un6_0_0_axb_39),.CI(un6_0_0_cry_38),.O(un6_0_0_s_39));
  MUXCY_L un6_0_0_cry_39_cZ(.DI(un6_0_8[39:39]),.CI(un6_0_0_cry_38),.S(un6_0_0_axb_39),.LO(un6_0_0_cry_39));
  XORCY un6_0_0_s_38_cZ(.LI(un6_0_0_axb_38),.CI(un6_0_0_cry_37),.O(un6_0_0_s_38));
  MUXCY_L un6_0_0_cry_38_cZ(.DI(un6_0_0_o5_37),.CI(un6_0_0_cry_37),.S(un6_0_0_axb_38),.LO(un6_0_0_cry_38));
  XORCY un6_0_0_s_37_cZ(.LI(un6_0_0_axb_37),.CI(un6_0_0_cry_36),.O(un6_0_0_s_37));
  MUXCY_L un6_0_0_cry_37_cZ(.DI(un6_0_9_s_21_RNIM4BU_O5),.CI(un6_0_0_cry_36),.S(un6_0_0_axb_37),.LO(un6_0_0_cry_37));
  XORCY un6_0_0_s_36_cZ(.LI(un6_0_0_axb_36),.CI(un6_0_0_cry_35),.O(un6_0_0_s_36));
  MUXCY_L un6_0_0_cry_36_cZ(.DI(un6_0_0_cry_36_RNO),.CI(un6_0_0_cry_35),.S(un6_0_0_axb_36),.LO(un6_0_0_cry_36));
  XORCY un6_0_0_s_35_cZ(.LI(un6_0_0_axb_35),.CI(un6_0_0_cry_34),.O(un6_0_0_s_35));
  MUXCY_L un6_0_0_cry_35_cZ(.DI(un6_0_0_cry_35_RNO),.CI(un6_0_0_cry_34),.S(un6_0_0_axb_35),.LO(un6_0_0_cry_35));
  XORCY un6_0_0_s_34_cZ(.LI(un6_0_0_axb_34),.CI(un6_0_0_cry_33),.O(un6_0_0_s_34));
  MUXCY_L un6_0_0_cry_34_cZ(.DI(un6_0_0_cry_34_RNO),.CI(un6_0_0_cry_33),.S(un6_0_0_axb_34),.LO(un6_0_0_cry_34));
  XORCY un6_0_0_s_33_cZ(.LI(un6_0_0_axb_33),.CI(un6_0_0_cry_32),.O(un6_0_0_s_33));
  MUXCY_L un6_0_0_cry_33_cZ(.DI(un6_0_0_cry_33_RNO),.CI(un6_0_0_cry_32),.S(un6_0_0_axb_33),.LO(un6_0_0_cry_33));
  XORCY un6_0_0_s_32_cZ(.LI(un6_0_0_axb_32),.CI(un6_0_0_cry_31),.O(un6_0_0_s_32));
  MUXCY_L un6_0_0_cry_32_cZ(.DI(un6_0_0_cry_32_RNO),.CI(un6_0_0_cry_31),.S(un6_0_0_axb_32),.LO(un6_0_0_cry_32));
  XORCY un6_0_0_s_31_cZ(.LI(un6_0_0_axb_31),.CI(un6_0_0_cry_30),.O(un6_0_0_s_31));
  MUXCY_L un6_0_0_cry_31_cZ(.DI(un6_0_0_cry_31_RNO),.CI(un6_0_0_cry_30),.S(un6_0_0_axb_31),.LO(un6_0_0_cry_31));
  XORCY un6_0_0_s_30_cZ(.LI(un6_0_0_axb_30),.CI(un6_0_0_cry_29),.O(un6_0_0_s_30));
  MUXCY_L un6_0_0_cry_30_cZ(.DI(un6_0_0_cry_30_RNO),.CI(un6_0_0_cry_29),.S(un6_0_0_axb_30),.LO(un6_0_0_cry_30));
  XORCY un6_0_0_s_29_cZ(.LI(un6_0_0_axb_29),.CI(un6_0_0_cry_28),.O(un6_0_0_s_29));
  MUXCY_L un6_0_0_cry_29_cZ(.DI(un6_0_0_cry_29_RNO),.CI(un6_0_0_cry_28),.S(un6_0_0_axb_29),.LO(un6_0_0_cry_29));
  XORCY un6_0_0_s_28_cZ(.LI(un6_0_0_axb_28),.CI(un6_0_0_cry_27),.O(un6_0_0_s_28));
  MUXCY_L un6_0_0_cry_28_cZ(.DI(un6_0_0_o5_27),.CI(un6_0_0_cry_27),.S(un6_0_0_axb_28),.LO(un6_0_0_cry_28));
  MUXCY_L un6_0_0_cry_27_cZ(.DI(un6_0_0_o5_26),.CI(un6_0_0_cry_26),.S(un6_0_0_axb_27),.LO(un6_0_0_cry_27));
  MUXCY_L un6_0_0_cry_26_cZ(.DI(un6_0_0_o5_25),.CI(un6_0_0_cry_25),.S(un6_0_0_axb_26),.LO(un6_0_0_cry_26));
  MUXCY_L un6_0_0_cry_25_cZ(.DI(un6_0_0_o5_24),.CI(un6_0_0_cry_24),.S(un6_0_0_axb_25),.LO(un6_0_0_cry_25));
  MUXCY_L un6_0_0_cry_24_cZ(.DI(un6_0_0_o5_23),.CI(un6_0_0_cry_23),.S(un6_0_0_axb_24),.LO(un6_0_0_cry_24));
  MUXCY_L un6_0_0_cry_23_cZ(.DI(un6_0_0_o5_22),.CI(un6_0_0_cry_22),.S(un6_0_0_axb_23),.LO(un6_0_0_cry_23));
  MUXCY_L un6_0_0_cry_22_cZ(.DI(un6_0_0_o5_21),.CI(un6_0_0_cry_21),.S(un6_0_0_axb_22),.LO(un6_0_0_cry_22));
  MUXCY_L un6_0_0_cry_21_cZ(.DI(un6_0_0_o5_20),.CI(un6_0_0_cry_20),.S(un6_0_0_axb_21),.LO(un6_0_0_cry_21));
  MUXCY_L un6_0_0_cry_20_cZ(.DI(un6_0_0_o5_19),.CI(un6_0_0_cry_19),.S(un6_0_0_axb_20),.LO(un6_0_0_cry_20));
  MUXCY_L un6_0_0_cry_19_cZ(.DI(un6_0_0_o5_18),.CI(un6_0_0_cry_18),.S(un6_0_0_axb_19),.LO(un6_0_0_cry_19));
  MUXCY_L un6_0_0_cry_18_cZ(.DI(un6_0_0_o5_17),.CI(un6_0_0_cry_17),.S(un6_0_0_axb_18),.LO(un6_0_0_cry_18));
  MUXCY_L un6_0_0_cry_17_cZ(.DI(un6_0_0_o5_16),.CI(un6_0_0_cry_16),.S(un6_0_0_axb_17),.LO(un6_0_0_cry_17));
  MUXCY_L un6_0_0_cry_16_cZ(.DI(un6_0_0_o5_15),.CI(un6_0_0_cry_15),.S(un6_0_0_axb_16),.LO(un6_0_0_cry_16));
  MUXCY_L un6_0_0_cry_15_cZ(.DI(un6_0_0_o5_14),.CI(un6_0_0_cry_14),.S(un6_0_0_axb_15),.LO(un6_0_0_cry_15));
  MUXCY_L un6_0_0_cry_14_cZ(.DI(un6_0_0_o5_13),.CI(un6_0_0_cry_13),.S(un6_0_0_axb_14),.LO(un6_0_0_cry_14));
  MUXCY_L un6_0_0_cry_13_cZ(.DI(un6_0_0_o5_12),.CI(un6_0_0_cry_12),.S(un6_0_0_axb_13),.LO(un6_0_0_cry_13));
  MUXCY_L un6_0_0_cry_12_cZ(.DI(un6_0_0_axb_11_lut6_2_O5),.CI(un6_0_0_cry_11),.S(un6_0_0_axb_12),.LO(un6_0_0_cry_12));
  MUXCY_L un6_0_0_cry_11_cZ(.DI(GND),.CI(un6_0_0_cry_10),.S(un6_0_0_axb_11),.LO(un6_0_0_cry_11));
  MUXCY_L un6_0_0_cry_10_cZ(.DI(un6_0_6[10:10]),.CI(un6_0_0_cry_9),.S(un6_0_0_axb_10),.LO(un6_0_0_cry_10));
  MUXCY_L un6_0_0_cry_9_cZ(.DI(un6_0_6[9:9]),.CI(un6_0_0_cry_8),.S(un6_0_0_axb_9),.LO(un6_0_0_cry_9));
  MUXCY_L un6_0_0_cry_8_cZ(.DI(un6_0_6[8:8]),.CI(un6_0_0_cry_7),.S(un6_0_0_axb_8),.LO(un6_0_0_cry_8));
  MUXCY_L un6_0_0_cry_7_cZ(.DI(un6_0_6[7:7]),.CI(un6_0_0_cry_6),.S(un6_0_0_axb_7),.LO(un6_0_0_cry_7));
  MUXCY_L un6_0_0_cry_6_cZ(.DI(GND),.CI(un6_0_0_cry_5),.S(un6_0_0_cry_6_sf),.LO(un6_0_0_cry_6));
  MUXCY_L un6_0_0_cry_5_cZ(.DI(GND),.CI(un6_0_0_cry_4),.S(un6_0_6[5:5]),.LO(un6_0_0_cry_5));
  MUXCY_L un6_0_0_cry_4_cZ(.DI(GND),.CI(un6_0_0_cry_3),.S(N_2381_i),.LO(un6_0_0_cry_4));
  MUXCY_L un6_0_0_cry_3_cZ(.DI(GND),.CI(un6_0_0_cry_2),.S(N_2384_i),.LO(un6_0_0_cry_3));
  MUXCY_L un6_0_0_cry_2_cZ(.DI(GND),.CI(un6_0_0_cry_1),.S(N_2387_i),.LO(un6_0_0_cry_2));
  MUXCY_L un6_0_0_cry_1_cZ(.DI(GND),.CI(un6_0_0_cry_0),.S(N_2390_i),.LO(un6_0_0_cry_1));
  MUXCY_L un6_0_0_cry_0_cZ(.DI(GND),.CI(VCC),.S(N_2393_i),.LO(un6_0_0_cry_0));
  XORCY un7_0_10_s_27(.LI(un7_0_10_s_27_true),.CI(un7_0_10_cry_26),.O(un7_0_10[45:45]));
  XORCY un7_0_10_s_26(.LI(un7_0_10_axb_26),.CI(un7_0_10_cry_25),.O(un7_0_10[44:44]));
  MUXCY_L un7_0_10_cry_26_cZ(.DI(GND),.CI(un7_0_10_cry_25),.S(un7_0_10_axb_26),.LO(un7_0_10_cry_26));
  XORCY un7_0_10_s_25(.LI(N_3385_i),.CI(un7_0_10_cry_24),.O(un7_0_10[43:43]));
  MUXCY_L un7_0_10_cry_25_cZ(.DI(VCC),.CI(un7_0_10_cry_24),.S(N_3385_i),.LO(un7_0_10_cry_25));
  XORCY un7_0_10_s_24(.LI(N_3387_i),.CI(un7_0_10_cry_23),.O(un7_0_10[42:42]));
  MUXCY_L un7_0_10_cry_24_cZ(.DI(VCC),.CI(un7_0_10_cry_23),.S(N_3387_i),.LO(un7_0_10_cry_24));
  XORCY un7_0_10_s_23(.LI(un7_0_10_axb_23),.CI(un7_0_10_cry_22),.O(un7_0_10[41:41]));
  MUXCY_L un7_0_10_cry_23_cZ(.DI(ZFF_X1[13:13]),.CI(un7_0_10_cry_22),.S(un7_0_10_axb_23),.LO(un7_0_10_cry_23));
  XORCY un7_0_10_s_22(.LI(un7_0_10_axb_22),.CI(un7_0_10_cry_21),.O(un7_0_10[40:40]));
  MUXCY_L un7_0_10_cry_22_cZ(.DI(un7_0_10_o5_21),.CI(un7_0_10_cry_21),.S(un7_0_10_axb_22),.LO(un7_0_10_cry_22));
  XORCY un7_0_10_s_21(.LI(un7_0_10_axb_21),.CI(un7_0_10_cry_20),.O(un7_0_10[39:39]));
  MUXCY_L un7_0_10_cry_21_cZ(.DI(un7_0_10_o5_20),.CI(un7_0_10_cry_20),.S(un7_0_10_axb_21),.LO(un7_0_10_cry_21));
  XORCY un7_0_10_s_20(.LI(un7_0_10_axb_20),.CI(un7_0_10_cry_19),.O(un7_0_10[38:38]));
  MUXCY_L un7_0_10_cry_20_cZ(.DI(un7_0_10_o5_19),.CI(un7_0_10_cry_19),.S(un7_0_10_axb_20),.LO(un7_0_10_cry_20));
  XORCY un7_0_10_s_19(.LI(un7_0_10_axb_19),.CI(un7_0_10_cry_18),.O(un7_0_10[37:37]));
  MUXCY_L un7_0_10_cry_19_cZ(.DI(un7_0_10_o5_18),.CI(un7_0_10_cry_18),.S(un7_0_10_axb_19),.LO(un7_0_10_cry_19));
  XORCY un7_0_10_s_18(.LI(un7_0_10_axb_18),.CI(un7_0_10_cry_17),.O(un7_0_10[36:36]));
  MUXCY_L un7_0_10_cry_18_cZ(.DI(un7_0_10_o5_17),.CI(un7_0_10_cry_17),.S(un7_0_10_axb_18),.LO(un7_0_10_cry_18));
  XORCY un7_0_10_s_17(.LI(un7_0_10_axb_17),.CI(un7_0_10_cry_16),.O(un7_0_10[35:35]));
  MUXCY_L un7_0_10_cry_17_cZ(.DI(un7_0_10_o5_16),.CI(un7_0_10_cry_16),.S(un7_0_10_axb_17),.LO(un7_0_10_cry_17));
  XORCY un7_0_10_s_16(.LI(un7_0_10_axb_16),.CI(un7_0_10_cry_15),.O(un7_0_10[34:34]));
  MUXCY_L un7_0_10_cry_16_cZ(.DI(un7_0_10_o5_15),.CI(un7_0_10_cry_15),.S(un7_0_10_axb_16),.LO(un7_0_10_cry_16));
  XORCY un7_0_10_s_15(.LI(un7_0_10_axb_15),.CI(un7_0_10_cry_14),.O(un7_0_10[33:33]));
  MUXCY_L un7_0_10_cry_15_cZ(.DI(un7_0_10_o5_14),.CI(un7_0_10_cry_14),.S(un7_0_10_axb_15),.LO(un7_0_10_cry_15));
  XORCY un7_0_10_s_14(.LI(un7_0_10_axb_14),.CI(un7_0_10_cry_13),.O(un7_0_10[32:32]));
  MUXCY_L un7_0_10_cry_14_cZ(.DI(un7_0_10_cry_14_RNO),.CI(un7_0_10_cry_13),.S(un7_0_10_axb_14),.LO(un7_0_10_cry_14));
  XORCY un7_0_10_s_13(.LI(un7_0_10_axb_13),.CI(un7_0_10_cry_12),.O(un7_0_10[31:31]));
  MUXCY_L un7_0_10_cry_13_cZ(.DI(un7_0_10_cry_13_RNO),.CI(un7_0_10_cry_12),.S(un7_0_10_axb_13),.LO(un7_0_10_cry_13));
  XORCY un7_0_10_s_12(.LI(un7_0_10_axb_12),.CI(un7_0_10_cry_11),.O(un7_0_10[30:30]));
  MUXCY_L un7_0_10_cry_12_cZ(.DI(un7_0_10_cry_12_RNO),.CI(un7_0_10_cry_11),.S(un7_0_10_axb_12),.LO(un7_0_10_cry_12));
  XORCY un7_0_10_s_11(.LI(un7_0_10_axb_11),.CI(un7_0_10_cry_10),.O(un7_0_10[29:29]));
  MUXCY_L un7_0_10_cry_11_cZ(.DI(N_2197_i),.CI(un7_0_10_cry_10),.S(un7_0_10_axb_11),.LO(un7_0_10_cry_11));
  XORCY un7_0_10_s_10(.LI(un7_0_10_axb_10),.CI(un7_0_10_cry_9),.O(un7_0_10[28:28]));
  MUXCY_L un7_0_10_cry_10_cZ(.DI(ZFF_X1[0:0]),.CI(un7_0_10_cry_9),.S(un7_0_10_axb_10),.LO(un7_0_10_cry_10));
  XORCY un7_0_10_s_9(.LI(un7_0_10_axb_9),.CI(un7_0_10_cry_8),.O(un7_0_10[27:27]));
  MUXCY_L un7_0_10_cry_9_cZ(.DI(GND),.CI(un7_0_10_cry_8),.S(un7_0_10_axb_9),.LO(un7_0_10_cry_9));
  XORCY un7_0_10_s_8(.LI(un7_0_10_axb_8),.CI(un7_0_10_cry_7),.O(un7_0_10[26:26]));
  MUXCY_L un7_0_10_cry_8_cZ(.DI(GND),.CI(un7_0_10_cry_7),.S(un7_0_10_axb_8),.LO(un7_0_10_cry_8));
  XORCY un7_0_10_s_7(.LI(un7_0_10_axb_7),.CI(un7_0_10_cry_6),.O(un7_0_10[25:25]));
  MUXCY_L un7_0_10_cry_7_cZ(.DI(GND),.CI(un7_0_10_cry_6),.S(un7_0_10_axb_7),.LO(un7_0_10_cry_7));
  XORCY un7_0_10_s_6(.LI(un7_0_10_axb_6),.CI(un7_0_10_cry_5),.O(un7_0_10[24:24]));
  MUXCY_L un7_0_10_cry_6_cZ(.DI(ZFF_X1[16:16]),.CI(un7_0_10_cry_5),.S(un7_0_10_axb_6),.LO(un7_0_10_cry_6));
  XORCY un7_0_10_s_5(.LI(un7_0_10_axb_5),.CI(un7_0_10_cry_4),.O(un7_0_10[23:23]));
  MUXCY_L un7_0_10_cry_5_cZ(.DI(ZFF_X1[16:16]),.CI(un7_0_10_cry_4),.S(un7_0_10_axb_5),.LO(un7_0_10_cry_5));
  XORCY un7_0_10_s_4(.LI(un7_0_10_axb_4),.CI(un7_0_10_cry_3),.O(un7_0_10[22:22]));
  MUXCY_L un7_0_10_cry_4_cZ(.DI(ZFF_X1[16:16]),.CI(un7_0_10_cry_3),.S(un7_0_10_axb_4),.LO(un7_0_10_cry_4));
  XORCY un7_0_10_s_3(.LI(un7_0_10_axb_3),.CI(un7_0_10_cry_2),.O(un7_0_10[21:21]));
  MUXCY_L un7_0_10_cry_3_cZ(.DI(GND),.CI(un7_0_10_cry_2),.S(un7_0_10_axb_3),.LO(un7_0_10_cry_3));
  XORCY un7_0_10_s_2(.LI(un7_0_10_axb_2),.CI(un7_0_10_cry_1),.O(un7_0_10[20:20]));
  MUXCY_L un7_0_10_cry_2_cZ(.DI(GND),.CI(un7_0_10_cry_1),.S(un7_0_10_axb_2),.LO(un7_0_10_cry_2));
  XORCY un7_0_10_s_1(.LI(un7_0_10_axb_1),.CI(un7_0_10_cry_0),.O(un7_0_10[19:19]));
  MUXCY_L un7_0_10_cry_1_cZ(.DI(un7_0_10_cry_1_RNO),.CI(un7_0_10_cry_0),.S(un7_0_10_axb_1),.LO(un7_0_10_cry_1));
  MUXCY_L un7_0_10_cry_0_cZ(.DI(un7_0_10_cry_0_RNO),.CI(GND),.S(un7_0_10[18:18]),.LO(un7_0_10_cry_0));
  BUFG state_reg_ret_5_cb_cZ(.I(un1_q_reg_2_c),.O(state_reg_ret_5_cb));
  LUT4 un10_axb_11_lut6_2_o6(.I0(ZFF_Y2[11:11]),.I1(un10_8[17:17]),.I2(un10_29),.I3(un10_6[17:17]),.O(un10_axb_11));
defparam un10_axb_11_lut6_2_o6.INIT=16'h9669;
  LUT3 un10_axb_11_lut6_2_o5(.I0(ZFF_Y2[11:11]),.I1(un10_8[17:17]),.I2(un10_29),.O(un10_axb_11_lut6_2_O5));
defparam un10_axb_11_lut6_2_o5.INIT=8'hD4;
  LUT2 un8_0_0_axb_11_lut6_2_o6(.I0(un8_0_8[11:11]),.I1(un8_0_6[11:11]),.O(un8_0_0_axb_11));
defparam un8_0_0_axb_11_lut6_2_o6.INIT=4'h6;
  LUT2 un8_0_0_axb_11_lut6_2_o5(.I0(un8_0_8[11:11]),.I1(un8_0_6[11:11]),.O(un8_0_0_axb_11_lut6_2_O5));
defparam un8_0_0_axb_11_lut6_2_o5.INIT=4'h8;
  LUT2 un6_0_0_axb_11_lut6_2_o6(.I0(un6_0_8[11:11]),.I1(un6_0_6[11:11]),.O(un6_0_0_axb_11));
defparam un6_0_0_axb_11_lut6_2_o6.INIT=4'h6;
  LUT2 un6_0_0_axb_11_lut6_2_o5(.I0(un6_0_8[11:11]),.I1(un6_0_6[11:11]),.O(un6_0_0_axb_11_lut6_2_O5));
defparam un6_0_0_axb_11_lut6_2_o5.INIT=4'h8;
  LUT4 un8_0_8_s_26_RNIUCD71_o6(.I0(un8_0_8[35:35]),.I1(un8_0_8[36:36]),.I2(un8_0_9[35:35]),.I3(un8_0_9[36:36]),.O(un8_0_0_axb_36));
defparam un8_0_8_s_26_RNIUCD71_o6.INIT=16'h6C93;
  LUT2 un8_0_8_s_26_RNIUCD71_o5(.I0(un8_0_8[36:36]),.I1(un8_0_9[36:36]),.O(un8_0_8_s_26_RNIUCD71_O5));
defparam un8_0_8_s_26_RNIUCD71_o5.INIT=4'hE;
  LUT4 un6_0_9_s_21_RNIM4BU_o6(.I0(un6_0_8[35:35]),.I1(un6_0_8[36:36]),.I2(un6_0_9[35:35]),.I3(un6_0_9[36:36]),.O(un6_0_0_axb_36));
defparam un6_0_9_s_21_RNIM4BU_o6.INIT=16'h6C93;
  LUT2 un6_0_9_s_21_RNIM4BU_o5(.I0(un6_0_8[36:36]),.I1(un6_0_9[36:36]),.O(un6_0_9_s_21_RNIM4BU_O5));
defparam un6_0_9_s_21_RNIM4BU_o5.INIT=4'hE;
  LUT4 un9_axb_1_lut6_2_o6(.I0(un9_8[6:6]),.I1(ZFF_Y1[3:3]),.I2(un9_8[7:7]),.I3(un9_10[8:8]),.O(un9_axb_1));
defparam un9_axb_1_lut6_2_o6.INIT=16'h6669;
  LUT3 un9_axb_1_lut6_2_o5(.I0(ZFF_Y1[3:3]),.I1(un9_8[7:7]),.I2(un9_10[8:8]),.O(un9_6[3:3]));
defparam un9_axb_1_lut6_2_o5.INIT=8'h56;
  LUT4 un9_axb_2_lut6_2_o6(.I0(ZFF_Y1[4:4]),.I1(ZFF_Y1[3:3]),.I2(un9_8[7:7]),.I3(un9_10[8:8]),.O(un9_axb_2));
defparam un9_axb_2_lut6_2_o6.INIT=16'h5A59;
  LUT4 un9_axb_2_lut6_2_o5(.I0(ZFF_Y1[4:4]),.I1(ZFF_Y1[3:3]),.I2(un9_8[7:7]),.I3(un9_10[8:8]),.O(un9_6[4:4]));
defparam un9_axb_2_lut6_2_o5.INIT=16'h5556;
  LUT3 un7_0_0_axb_10_lut6_2_o6(.I0(ZFF_X1[1:1]),.I1(un7_0_6[10:10]),.I2(un7_0_8[10:10]),.O(un7_0_0_axb_10));
defparam un7_0_0_axb_10_lut6_2_o6.INIT=8'h96;
  LUT3 un7_0_0_axb_10_lut6_2_o5(.I0(ZFF_X1[1:1]),.I1(un7_0_6[10:10]),.I2(un7_0_8[10:10]),.O(un7_0_0_axb_10_lut6_2_O5));
defparam un7_0_0_axb_10_lut6_2_o5.INIT=8'hE8;
  LUT5 sum_stg_a_lut6_2_o6(.I0(q_reg_i_1[0:0]),.I1(q_reg[2:2]),.I2(q_reg_i_1[1:1]),.I3(q_reg_i_1[2:2]),.I4(state_reg),.O(sum_stg_a));
defparam sum_stg_a_lut6_2_o6.INIT=32'hCC800000;
  LUT3 sum_stg_a_lut6_2_o5(.I0(q_reg_i_1[1:1]),.I1(q_reg_i_1[2:2]),.I2(state_reg),.O(filter_done));
defparam sum_stg_a_lut6_2_o5.INIT=8'h10;
  LUT4 trunc_out_lut6_2_o6(.I0(q_reg_i_1[0:0]),.I1(q_reg_i_1[1:1]),.I2(q_reg_i_1[2:2]),.I3(state_reg),.O(trunc_out));
defparam trunc_out_lut6_2_o6.INIT=16'h0400;
  LUT3 trunc_out_lut6_2_o5(.I0(state_reg_ret_4),.I1(q_reg_i_1[2:2]),.I2(state_reg),.O(trunc_prods));
defparam trunc_out_lut6_2_o5.INIT=8'h40;
  LUT4 desc498(.I0(q_reg[0:0]),.I1(q_reg_i_1[1:1]),.I2(q_reg_i_1[2:2]),.I3(state_reg),.O(q_next[0:0]));
defparam desc498.INIT=16'h54AA;
  LUT5 desc499(.I0(q_reg[1:1]),.I1(q_reg[0:0]),.I2(q_reg_i_1[1:1]),.I3(q_reg_i_1[2:2]),.I4(state_reg),.O(q_next[1:1]));
defparam desc499.INIT=32'h6660AAAA;
  LUT5 desc500(.I0(q_reg[1:1]),.I1(q_reg[0:0]),.I2(q_reg_i_1[1:1]),.I3(q_reg_i_1[2:2]),.I4(state_reg),.O(q_next_i[1:1]));
defparam desc500.INIT=32'h999F5555;
  LUT4 desc501(.I0(q_reg[0:0]),.I1(q_reg_i_1[1:1]),.I2(q_reg_i_1[2:2]),.I3(state_reg),.O(q_next_i[0:0]));
defparam desc501.INIT=16'hAB55;
  LUT5 un9_axb_3_lut6_2_o6(.I0(ZFF_Y1[5:5]),.I1(ZFF_Y1[4:4]),.I2(ZFF_Y1[3:3]),.I3(un9_8[7:7]),.I4(un9_10[8:8]),.O(un9_axb_3));
defparam un9_axb_3_lut6_2_o6.INIT=32'hA5A55A59;
  LUT5 un9_axb_3_lut6_2_o5(.I0(ZFF_Y1[5:5]),.I1(ZFF_Y1[4:4]),.I2(ZFF_Y1[3:3]),.I3(un9_8[7:7]),.I4(un9_10[8:8]),.O(un9_6[5:5]));
defparam un9_axb_3_lut6_2_o5.INIT=32'hAAAA5556;
  LUT2 desc502(.I0(ZFF_Y2[6:6]),.I1(ZFF_Y2[0:0]),.O(un10_6_i[6:6]));
defparam desc502.INIT=4'h6;
  LUT2 desc503(.I0(ZFF_Y2[6:6]),.I1(ZFF_Y2[0:0]),.O(un10_6[6:6]));
defparam desc503.INIT=4'h9;
  LUT4 desc504(.I0(ZFF_Y2[7:7]),.I1(ZFF_Y2[6:6]),.I2(ZFF_Y2[0:0]),.I3(ZFF_Y2[1:1]),.O(un10_axb_1));
defparam desc504.INIT=16'hA659;
  LUT2 desc505(.I0(ZFF_Y2[6:6]),.I1(ZFF_Y2[0:0]),.O(un10_6[7:7]));
defparam desc505.INIT=4'h2;
  LUT5 desc506(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[7:7]),.I2(ZFF_Y2[0:0]),.I3(ZFF_Y2[2:2]),.I4(ZFF_Y2[1:1]),.O(un10_axb_2));
defparam desc506.INIT=32'h5AA59669;
  LUT3 desc507(.I0(ZFF_Y2[8:8]),.I1(ZFF_Y2[0:0]),.I2(ZFF_Y2[2:2]),.O(un10_6[8:8]));
defparam desc507.INIT=8'h96;
endmodule