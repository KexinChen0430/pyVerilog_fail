module.ids[id]))
    */
   /*metav_generated:*/
   assign ignored = "This code is ignored by the lexer";
   syntax errors are ignored;
   Lexer errors are also ignored: ¤;
   /*:metav_generated*/
endmodule