module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_aa
		ent_aa inst_aa (
		);
		// End of Generated Instance Port Map for inst_aa
		// Generated Instance Port Map for inst_ab
		ent_ab inst_ab (
		);
		// End of Generated Instance Port Map for inst_ab
		// Generated Instance Port Map for inst_ac
		ent_ac inst_ac (
		);
		// End of Generated Instance Port Map for inst_ac
		// Generated Instance Port Map for inst_ad
		ent_ad inst_ad (
		);
		// End of Generated Instance Port Map for inst_ad
		// Generated Instance Port Map for inst_ae
		ent_ae inst_ae (
		);
		// End of Generated Instance Port Map for inst_ae
endmodule