module outputs
  wire [127 : 0] wmemiM_MData;
  wire [35 : 0] wmemiM_MAddr;
  wire [31 : 0] wci_s_0_SData,
		wci_s_1_SData,
		wci_s_2_SData,
		wci_s_3_SData,
		wci_s_4_SData,
		wci_s_5_SData,
		wci_s_6_SData,
		wci_s_7_SData,
		wmiM0_MData,
		wmiM0_MFlag,
		wmiM1_MData,
		wmiM1_MFlag,
		wsi_m_dac_MData;
  wire [15 : 0] wmemiM_MDataByteEn;
  wire [13 : 0] wmiM0_MAddr, wmiM1_MAddr;
  wire [11 : 0] wmemiM_MBurstLength,
		wmiM0_MBurstLength,
		wmiM1_MBurstLength,
		wsi_m_dac_MBurstLength;
  wire [7 : 0] wsi_m_dac_MReqInfo;
  wire [3 : 0] wmiM0_MDataByteEn, wmiM1_MDataByteEn, wsi_m_dac_MByteEn;
  wire [2 : 0] wmemiM_MCmd, wmiM0_MCmd, wmiM1_MCmd, wsi_m_dac_MCmd;
  wire [1 : 0] wci_s_0_SFlag,
	       wci_s_0_SResp,
	       wci_s_1_SFlag,
	       wci_s_1_SResp,
	       wci_s_2_SFlag,
	       wci_s_2_SResp,
	       wci_s_3_SFlag,
	       wci_s_3_SResp,
	       wci_s_4_SFlag,
	       wci_s_4_SResp,
	       wci_s_5_SFlag,
	       wci_s_5_SResp,
	       wci_s_6_SFlag,
	       wci_s_6_SResp,
	       wci_s_7_SFlag,
	       wci_s_7_SResp;
  wire wci_s_0_SThreadBusy,
       wci_s_1_SThreadBusy,
       wci_s_2_SThreadBusy,
       wci_s_3_SThreadBusy,
       wci_s_4_SThreadBusy,
       wci_s_5_SThreadBusy,
       wci_s_6_SThreadBusy,
       wci_s_7_SThreadBusy,
       wmemiM_MDataLast,
       wmemiM_MDataValid,
       wmemiM_MReqLast,
       wmemiM_MReset_n,
       wmiM0_MAddrSpace,
       wmiM0_MDataLast,
       wmiM0_MDataValid,
       wmiM0_MReqInfo,
       wmiM0_MReqLast,
       wmiM0_MReset_n,
       wmiM1_MAddrSpace,
       wmiM1_MDataLast,
       wmiM1_MDataValid,
       wmiM1_MReqInfo,
       wmiM1_MReqLast,
       wmiM1_MReset_n,
       wsi_m_dac_MBurstPrecise,
       wsi_m_dac_MReqLast,
       wsi_m_dac_MReset_n,
       wsi_s_adc_SReset_n,
       wsi_s_adc_SThreadBusy;
  // Instantiate the wip-compliant app
  ocpi_app #(.hasDebugLogic(hasDebugLogic)) app(
				      .wci0_MReset_n(RST_N_rst_2),
				      .wci1_MReset_n(RST_N_rst_3),
				      .wci2_MReset_n(RST_N_rst_4),
				      .wci3_MReset_n(RST_N_rst_5),
				      .wci4_MReset_n(RST_N_rst_6),
				      .wci5_MReset_n(RST_N_rst_7),
				      .wci_Clk(CLK),
				      .wci0_MAddr(wci_s_2_MAddr),
				      .wci0_MAddrSpace(wci_s_2_MAddrSpace),
				      .wci0_MByteEn(wci_s_2_MByteEn),
				      .wci0_MCmd(wci_s_2_MCmd),
				      .wci0_MData(wci_s_2_MData),
				      .wci0_MFlag(wci_s_2_MFlag),
				      .wci1_MAddr(wci_s_3_MAddr),
				      .wci1_MAddrSpace(wci_s_3_MAddrSpace),
				      .wci1_MByteEn(wci_s_3_MByteEn),
				      .wci1_MCmd(wci_s_3_MCmd),
				      .wci1_MData(wci_s_3_MData),
				      .wci1_MFlag(wci_s_3_MFlag),
				      .wci2_MAddr(wci_s_4_MAddr),
				      .wci2_MAddrSpace(wci_s_4_MAddrSpace),
				      .wci2_MByteEn(wci_s_4_MByteEn),
				      .wci2_MCmd(wci_s_4_MCmd),
				      .wci2_MData(wci_s_4_MData),
				      .wci2_MFlag(wci_s_4_MFlag),
				      .wci3_MAddr(wci_s_5_MAddr),
				      .wci3_MAddrSpace(wci_s_5_MAddrSpace),
				      .wci3_MByteEn(wci_s_5_MByteEn),
				      .wci3_MCmd(wci_s_5_MCmd),
				      .wci3_MData(wci_s_5_MData),
				      .wci3_MFlag(wci_s_5_MFlag),
				      .wci4_MAddr(wci_s_6_MAddr),
				      .wci4_MAddrSpace(wci_s_6_MAddrSpace),
				      .wci4_MByteEn(wci_s_6_MByteEn),
				      .wci4_MCmd(wci_s_6_MCmd),
				      .wci4_MData(wci_s_6_MData),
				      .wci4_MFlag(wci_s_6_MFlag),
				      .wci5_MAddr(wci_s_7_MAddr),
				      .wci5_MAddrSpace(wci_s_7_MAddrSpace),
				      .wci5_MByteEn(wci_s_7_MByteEn),
				      .wci5_MCmd(wci_s_7_MCmd),
				      .wci5_MData(wci_s_7_MData),
				      .wci5_MFlag(wci_s_7_MFlag),
				      .wmemi0_SData(wmemiM_SData),
				      .wmemi0_SResp(wmemiM_SResp),
				      .wmiM0_SData(wmiM0_SData),
				      .wmiM0_SFlag(wmiM0_SFlag),
				      .wmiM0_SResp(wmiM0_SResp),
				      .wmiM1_SData(wmiM1_SData),
				      .wmiM1_SFlag(wmiM1_SFlag),
				      .wmiM1_SResp(wmiM1_SResp),
				      .adc_MBurstLength(wsi_s_adc_MBurstLength),
				      .adc_MByteEn(wsi_s_adc_MByteEn),
				      .adc_MCmd(wsi_s_adc_MCmd),
				      .adc_MData(wsi_s_adc_MData),
				      .adc_MReqInfo(wsi_s_adc_MReqInfo),
				      .wmiM0_SThreadBusy(wmiM0_SThreadBusy),
				      .wmiM0_SDataThreadBusy(wmiM0_SDataThreadBusy),
				      .wmiM0_SRespLast(wmiM0_SRespLast),
				      .wmiM0_SReset_n(wmiM0_SReset_n),
				      .wmiM1_SThreadBusy(wmiM1_SThreadBusy),
				      .wmiM1_SDataThreadBusy(wmiM1_SDataThreadBusy),
				      .wmiM1_SRespLast(wmiM1_SRespLast),
				      .wmiM1_SReset_n(wmiM1_SReset_n),
				      .wmemi0_SRespLast(wmemiM_SRespLast),
				      .wmemi0_SCmdAccept(wmemiM_SCmdAccept),
				      .wmemi0_SDataAccept(wmemiM_SDataAccept),
				      .adc_MReqLast(wsi_s_adc_MReqLast),
				      .adc_MBurstPrecise(wsi_s_adc_MBurstPrecise),
				      .adc_MReset_n(wsi_s_adc_MReset_n),
				      .dac_SThreadBusy(wsi_m_dac_SThreadBusy),
				      .dac_SReset_n(wsi_m_dac_SReset_n),
				      .wci0_SResp(wci_s_2_SResp),
				      .wci0_SData(wci_s_2_SData),
				      .wci0_SThreadBusy(wci_s_2_SThreadBusy),
				      .wci0_SFlag(wci_s_2_SFlag),
				      .wci1_SResp(wci_s_3_SResp),
				      .wci1_SData(wci_s_3_SData),
				      .wci1_SThreadBusy(wci_s_3_SThreadBusy),
				      .wci1_SFlag(wci_s_3_SFlag),
				      .wci2_SResp(wci_s_4_SResp),
				      .wci2_SData(wci_s_4_SData),
				      .wci2_SThreadBusy(wci_s_4_SThreadBusy),
				      .wci2_SFlag(wci_s_4_SFlag),
				      .wci3_SResp(wci_s_5_SResp),
				      .wci3_SData(wci_s_5_SData),
				      .wci3_SThreadBusy(wci_s_5_SThreadBusy),
				      .wci3_SFlag(wci_s_5_SFlag),
				      .wci4_SResp(wci_s_6_SResp),
				      .wci4_SData(wci_s_6_SData),
				      .wci4_SThreadBusy(wci_s_6_SThreadBusy),
				      .wci4_SFlag(wci_s_6_SFlag),
				      .wci5_SResp(wci_s_7_SResp),
				      .wci5_SData(wci_s_7_SData),
				      .wci5_SThreadBusy(wci_s_7_SThreadBusy),
				      .wci5_SFlag(wci_s_7_SFlag),
				      .wmiM0_MCmd(wmiM0_MCmd),
				      .wmiM0_MReqLast(wmiM0_MReqLast),
				      .wmiM0_MReqInfo(wmiM0_MReqInfo),
				      .wmiM0_MAddrSpace(wmiM0_MAddrSpace),
				      .wmiM0_MAddr(wmiM0_MAddr),
				      .wmiM0_MBurstLength(wmiM0_MBurstLength),
				      .wmiM0_MDataValid(wmiM0_MDataValid),
				      .wmiM0_MDataLast(wmiM0_MDataLast),
				      .wmiM0_MData(wmiM0_MData),
				      .wmiM0_MDataByteEn(wmiM0_MDataByteEn),
				      .wmiM0_MFlag(wmiM0_MFlag),
				      .wmiM0_MReset_n(wmiM0_MReset_n),
				      .wmiM1_MCmd(wmiM1_MCmd),
				      .wmiM1_MReqLast(wmiM1_MReqLast),
				      .wmiM1_MReqInfo(wmiM1_MReqInfo),
				      .wmiM1_MAddrSpace(wmiM1_MAddrSpace),
				      .wmiM1_MAddr(wmiM1_MAddr),
				      .wmiM1_MBurstLength(wmiM1_MBurstLength),
				      .wmiM1_MDataValid(wmiM1_MDataValid),
				      .wmiM1_MDataLast(wmiM1_MDataLast),
				      .wmiM1_MData(wmiM1_MData),
				      .wmiM1_MDataByteEn(wmiM1_MDataByteEn),
				      .wmiM1_MFlag(wmiM1_MFlag),
				      .wmiM1_MReset_n(wmiM1_MReset_n),
				      .wmemi0_MCmd(wmemiM_MCmd),
				      .wmemi0_MReqLast(wmemiM_MReqLast),
				      .wmemi0_MAddr(wmemiM_MAddr),
				      .wmemi0_MBurstLength(wmemiM_MBurstLength),
				      .wmemi0_MDataValid(wmemiM_MDataValid),
				      .wmemi0_MDataLast(wmemiM_MDataLast),
				      .wmemi0_MData(wmemiM_MData),
				      .wmemi0_MDataByteEn(wmemiM_MDataByteEn),
				      .wmemi0_MReset_n(wmemiM_MReset_n),
				      .adc_SThreadBusy(wsi_s_adc_SThreadBusy),
				      .adc_SReset_n(wsi_s_adc_SReset_n),
				      .dac_MCmd(wsi_m_dac_MCmd),
				      .dac_MReqLast(wsi_m_dac_MReqLast),
				      .dac_MBurstPrecise(wsi_m_dac_MBurstPrecise),
				      .dac_MBurstLength(wsi_m_dac_MBurstLength),
				      .dac_MData(wsi_m_dac_MData),
				      .dac_MByteEn(wsi_m_dac_MByteEn),
				      .dac_MReqInfo(wsi_m_dac_MReqInfo),
				      .dac_MReset_n(wsi_m_dac_MReset_n));
endmodule