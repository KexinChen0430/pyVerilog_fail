module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for cgu_i
		cgu cgu_i (
		);
		// End of Generated Instance Port Map for cgu_i
		// Generated Instance Port Map for tmu_i
		tmu tmu_i (
		);
		// End of Generated Instance Port Map for tmu_i
endmodule