module ram_controller_phy_alt_mem_phy_mimic(
                         //Inputs
                         //Clocks
                         measure_clk,         // full rate clock from PLL
                         mimic_data_in,       // Input against which the VT variations
                                              // are tracked (e.g. memory clock)
                         // Active low reset
                         reset_measure_clk_n,
                         //Indicates that the mimic calibration sequence can start
                         seq_mmc_start,       // from sequencer
                         //Outputs
                         mmc_seq_done,        // mimic calibration finished for the current PLL phase
                         mmc_seq_value        // result value of the mimic calibration
        );
   input  wire measure_clk;
   input  wire mimic_data_in;
   input  wire reset_measure_clk_n;
   input  wire seq_mmc_start;
   output wire mmc_seq_done;
   output wire mmc_seq_value;
   function integer clogb2;
      input [31:0] value;
      for (clogb2=0; value>0; clogb2=clogb2+1)
          value = value >> 1;
   endfunction // clogb2
   // Parameters
   parameter NUM_MIMIC_SAMPLE_CYCLES = 6;
   parameter SHIFT_REG_COUNTER_WIDTH = clogb2(NUM_MIMIC_SAMPLE_CYCLES);
   reg [`MIMIC_FSM_WIDTH-1:0]           mimic_state;
   reg [2:0]                            seq_mmc_start_metastable;
   wire                                 start_edge_detected;
   (* altera_attribute=" -name fast_input_register OFF"*) reg [1:0] mimic_data_in_metastable;
   wire                                 mimic_data_in_sample;
   wire                                 shift_reg_data_out_all_ones;
   reg                                  mimic_done_out;
   reg                                  mimic_value_captured;
   reg [SHIFT_REG_COUNTER_WIDTH : 0]    shift_reg_counter;
   reg                                  shift_reg_enable;
   wire                                 shift_reg_data_in;
   reg                                  shift_reg_s_clr;
   wire                                 shift_reg_a_clr;
   reg [NUM_MIMIC_SAMPLE_CYCLES -1 : 0] shift_reg_data_out;
   // shift register which contains the sampled data
   always @(posedge measure_clk or posedge shift_reg_a_clr)
   begin
      if (shift_reg_a_clr == 1'b1)
      begin
          shift_reg_data_out    <= {NUM_MIMIC_SAMPLE_CYCLES{1'b0}};
      end
      else
      begin
         if (shift_reg_s_clr == 1'b1)
         begin
             shift_reg_data_out <= {NUM_MIMIC_SAMPLE_CYCLES{1'b0}};
         end
         else if (shift_reg_enable == 1'b1)
         begin
             shift_reg_data_out <= {(shift_reg_data_out[NUM_MIMIC_SAMPLE_CYCLES -2 : 0]), shift_reg_data_in};
         end
      end
   end
  // Metastable-harden mimic_start :
  always @(posedge measure_clk or negedge reset_measure_clk_n)
  begin
    if (reset_measure_clk_n == 1'b0)
    begin
        seq_mmc_start_metastable    <= 0;
    end
    else
    begin
        seq_mmc_start_metastable[0] <= seq_mmc_start;
        seq_mmc_start_metastable[1] <= seq_mmc_start_metastable[0];
        seq_mmc_start_metastable[2] <= seq_mmc_start_metastable[1];
    end
  end
  assign start_edge_detected =  seq_mmc_start_metastable[1]
                             && !seq_mmc_start_metastable[2];
  // Metastable-harden mimic_data_in :
  always @(posedge measure_clk or negedge reset_measure_clk_n)
  begin
    if (reset_measure_clk_n == 1'b0)
    begin
        mimic_data_in_metastable    <= 0;
    end
      //some mimic paths configurations have another flop inside the wysiwyg ioe
    else
    begin
        mimic_data_in_metastable[0] <= mimic_data_in;
        mimic_data_in_metastable[1] <= mimic_data_in_metastable[0];
    end
  end
  assign mimic_data_in_sample =  mimic_data_in_metastable[1];
  // Main FSM :
  always @(posedge measure_clk or negedge reset_measure_clk_n )
  begin
     if (reset_measure_clk_n == 1'b0)
     begin
         mimic_state           <= `MIMIC_IDLE;
         mimic_done_out        <= 1'b0;
         mimic_value_captured  <= 1'b0;
         shift_reg_counter     <= 0;
         shift_reg_enable      <= 1'b0;
         shift_reg_s_clr       <= 1'b0;
     end
     else
     begin
         case (mimic_state)
         `MIMIC_IDLE : begin
                           shift_reg_counter     <= 0;
                           mimic_done_out        <= 1'b0;
                           shift_reg_s_clr       <= 1'b1;
                           shift_reg_enable      <= 1'b1;
                           if (start_edge_detected == 1'b1)
                           begin
                               mimic_state       <= `MIMIC_SAMPLE;
                               shift_reg_counter <= shift_reg_counter + 1'b1;
                               shift_reg_s_clr   <= 1'b0;
                           end
                           else
                           begin
                               mimic_state <= `MIMIC_IDLE;
                           end
         end // case: MIMIC_IDLE
           `MIMIC_SAMPLE : begin
                               shift_reg_counter        <= shift_reg_counter + 1'b1;
                               if (shift_reg_counter == NUM_MIMIC_SAMPLE_CYCLES + 1)
                               begin
                                   mimic_done_out       <= 1'b1;
                                   mimic_value_captured <= shift_reg_data_out_all_ones; //captured only here
                                   shift_reg_enable     <= 1'b0;
                                   shift_reg_counter    <= shift_reg_counter;
                                   mimic_state          <= `MIMIC_SEND;
                               end
           end // case: MIMIC_SAMPLE
           `MIMIC_SEND : begin
                             mimic_done_out  <= 1'b1; //redundant statement, here just for readibility
                             mimic_state     <= `MIMIC_SEND1;
            /* mimic_value_captured will not change during MIMIC_SEND
               it will change next time mimic_done_out is asserted
               mimic_done_out will be reset during MIMIC_IDLE
               the purpose of the current state is to add one clock cycle
               mimic_done_out will be active for 2 measure_clk clock cycles, i.e
               the pulses duration will be just one sequencer clock cycle
               (which is half rate) */
           end // case: MIMIC_SEND
           // MIMIC_SEND1 and MIMIC_SEND2 extend the mimic_done_out signal by another 2 measure_clk_2x cycles
           // so it is a total of 4 measure clocks long (ie 2 half-rate clock cycles long in total)
           `MIMIC_SEND1 : begin
                              mimic_done_out  <= 1'b1; //redundant statement, here just for readibility
                              mimic_state     <= `MIMIC_SEND2;
           end
           `MIMIC_SEND2 : begin
                              mimic_done_out  <= 1'b1; //redundant statement, here just for readibility
                              mimic_state     <= `MIMIC_IDLE;
           end
           default : begin
                         mimic_state <= `MIMIC_IDLE;
           end
         endcase
     end
  end
  assign shift_reg_data_out_all_ones   = (( & shift_reg_data_out) == 1'b1) ? 1'b1
                                                                           : 1'b0;
  // Shift Register assignments
  assign shift_reg_data_in  =  mimic_data_in_sample;
  assign shift_reg_a_clr    =  !reset_measure_clk_n;
  // Output assignments
  assign mmc_seq_done    = mimic_done_out;
  assign mmc_seq_value   = mimic_value_captured;
endmodule