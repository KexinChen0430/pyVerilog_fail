module ks3e9b2 (
   input wire         sys_clk ,
   input wire         rst_n ,
   input wire [15:0]  ux36419 ,
   input wire         ep85b3b ,
   input wire         nt2d9dd ,
   input              fnd82ee ,
   output reg [31:0]  gof0cd8 ,
   output wire        zm866c1 ,
   output wire        ld6baf6        ) ;
reg              jc5d7b7 ;
reg              lqebdbb ;
reg              kd5eddb ;
reg [15:0]       vvf6edd ;
reg [15:0]       lsb76ee ;
reg [15:0]       ohbb773 ;
reg [31:0]       osdbb9d ;
reg [31:0]       blddce9 ;
reg [15:0]       viee74e ;
wire             ho73a72 ;
wire [31:0]      co9d392 ;
wire [15:0]      jpe9c91 ;
wire             qt4e48e ;
wire             go72475 ;
reg [15 : 0] ym923a9;
reg vx91d48;
reg xl8ea46;
reg ng1a6b;
reg ksa91b4;
reg by48da1;
reg [15 : 0] qg46d0b;
reg [15 : 0] an36858;
reg [15 : 0] anb42c4;
reg [31 : 0] ana1624;
reg [31 : 0] vkb125;
reg [15 : 0] vi5892b;
reg ykc495a;
reg [31 : 0] ou24ad1;
reg [15 : 0] zm25688;
reg mg2b443;
reg pf5a218;
reg [2047:0] necf6c2;
wire [16:0] ld7b613;
localparam qgdb09f = 17,nrd84f8 = 32'hfdffe42b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
assign ho73a72 = vx91d48 ;
always @(posedge sys_clk, negedge rst_n) begin   if (!rst_n) begin      jc5d7b7 <= 1'b0 ;      lqebdbb <= 1'b0 ;      kd5eddb <= 1'b0 ;   end   else  begin      jc5d7b7 <=  ykc495a ;      lqebdbb <=  jc5d7b7 ;      kd5eddb <=  ksa91b4 ;   end
end
always @(posedge sys_clk, negedge rst_n) begin   if (!rst_n)      vvf6edd <= 1'd0 ;   else if (ykc495a)      vvf6edd <= ym923a9 ;   else      vvf6edd <= qg46d0b ;
end
assign co9d392 = {qg46d0b, ym923a9} ;
always @* begin   blddce9 = ou24ad1 ;   osdbb9d = {vkb125[24],vkb125[25],vkb125[26],vkb125[27],vkb125[28],vkb125[29],vkb125[30],vkb125[31],        vkb125[16],vkb125[17],vkb125[18],vkb125[19],vkb125[20],vkb125[21],vkb125[22],vkb125[23],        vkb125[8],vkb125[9],vkb125[10],vkb125[11],vkb125[12],vkb125[13],vkb125[14],vkb125[15],        vkb125[0],vkb125[1],vkb125[2],vkb125[3],vkb125[4],vkb125[5],vkb125[6],vkb125[7] };   ohbb773 = 16'h32B9;   lsb76ee[0] = ana1624[31] ^ ana1624[29] ^ ana1624[28] ^ ana1624[26] ^ ana1624[23] ^ ana1624[21] ^ ana1624[20] ^               ana1624[15] ^ ana1624[13] ^ ana1624[12] ^ ana1624[8] ^ ana1624[4] ^ ana1624[0] ^ anb42c4[0] ;   lsb76ee[1] = ana1624[31] ^ ana1624[30] ^ ana1624[28] ^ ana1624[27] ^ ana1624[26] ^ ana1624[24] ^ ana1624[23] ^               ana1624[22] ^ ana1624[20] ^ ana1624[16] ^ ana1624[15] ^ ana1624[14] ^ ana1624[12] ^ ana1624[9] ^               ana1624[8] ^ ana1624[5] ^ ana1624[4] ^ ana1624[1] ^ ana1624[0] ^ anb42c4[1] ;   lsb76ee[2] = ana1624[31] ^ ana1624[29] ^ ana1624[28] ^ ana1624[27] ^ ana1624[25] ^ ana1624[24] ^ ana1624[23] ^               ana1624[21] ^ ana1624[17] ^ ana1624[16] ^ ana1624[15] ^ ana1624[13] ^ ana1624[10] ^ ana1624[9] ^               ana1624[6] ^ ana1624[5] ^ ana1624[2] ^ ana1624[1] ^ anb42c4[2] ;   lsb76ee[3] = ana1624[31] ^ ana1624[30] ^ ana1624[25] ^ ana1624[24] ^ ana1624[23] ^ ana1624[22] ^ ana1624[21] ^               ana1624[20] ^ ana1624[18] ^ ana1624[17] ^ ana1624[16] ^ ana1624[15] ^ ana1624[14] ^ ana1624[13] ^               ana1624[12] ^ ana1624[11] ^ ana1624[10] ^ ana1624[8] ^ ana1624[7] ^ ana1624[6] ^ ana1624[4] ^               ana1624[3] ^ ana1624[2] ^ ana1624[0] ^ anb42c4[3] ;   lsb76ee[4] = ana1624[31] ^ ana1624[26] ^ ana1624[25] ^ ana1624[24] ^ ana1624[23] ^ ana1624[22] ^ ana1624[21] ^               ana1624[19] ^ ana1624[18] ^ ana1624[17] ^ ana1624[16] ^ ana1624[15] ^ ana1624[14] ^ ana1624[13] ^               ana1624[12] ^ ana1624[11] ^ ana1624[9] ^ ana1624[8] ^ ana1624[7] ^ ana1624[5] ^ ana1624[4] ^               ana1624[3] ^ ana1624[1] ^ anb42c4[4] ;   lsb76ee[5] = ana1624[27] ^ ana1624[26] ^ ana1624[25] ^ ana1624[24] ^ ana1624[23] ^ ana1624[22] ^ ana1624[20] ^               ana1624[19] ^ ana1624[18] ^ ana1624[17] ^ ana1624[16] ^ ana1624[15] ^ ana1624[14] ^ ana1624[13] ^               ana1624[12] ^ ana1624[10] ^ ana1624[9] ^ ana1624[8] ^ ana1624[6] ^ ana1624[5] ^ ana1624[4] ^               ana1624[2] ^  anb42c4[5] ;   lsb76ee[6] = ana1624[28] ^ ana1624[27] ^ ana1624[26] ^ ana1624[25] ^ ana1624[24] ^ ana1624[23] ^ ana1624[21] ^               ana1624[20] ^ ana1624[19] ^ ana1624[18] ^ ana1624[17] ^ ana1624[16] ^ ana1624[15] ^ ana1624[14] ^               ana1624[13] ^ ana1624[11] ^ ana1624[10] ^ ana1624[9] ^ ana1624[7] ^ ana1624[6] ^ ana1624[5] ^               ana1624[3] ^ anb42c4[6] ;   lsb76ee[7] = ana1624[29] ^ ana1624[28] ^ ana1624[27] ^ ana1624[26] ^ ana1624[25] ^ ana1624[24] ^ ana1624[22] ^               ana1624[21] ^ ana1624[20] ^ ana1624[19] ^ ana1624[18] ^ ana1624[17] ^ ana1624[16] ^ ana1624[15] ^               ana1624[14] ^ ana1624[12] ^ ana1624[11] ^ ana1624[10] ^ ana1624[8] ^ ana1624[7] ^ ana1624[6] ^               ana1624[4] ^ anb42c4[7] ;   lsb76ee[8] = ana1624[30] ^ ana1624[29] ^ ana1624[28] ^ ana1624[27] ^ ana1624[26] ^ ana1624[25] ^ ana1624[23] ^               ana1624[22] ^ ana1624[21] ^ ana1624[20] ^ ana1624[19] ^ ana1624[18] ^ ana1624[17] ^ ana1624[16] ^               ana1624[15] ^ ana1624[13] ^ ana1624[12] ^ ana1624[11] ^ ana1624[9] ^ ana1624[8] ^ ana1624[7] ^               ana1624[5] ^ anb42c4[8] ;   lsb76ee[9] = ana1624[31] ^ ana1624[30] ^ ana1624[29] ^ ana1624[28] ^ ana1624[27] ^ ana1624[26] ^ ana1624[24] ^               ana1624[23] ^ ana1624[22] ^ ana1624[21] ^ ana1624[20] ^ ana1624[19] ^ ana1624[18] ^ ana1624[17] ^               ana1624[16] ^ ana1624[14] ^ ana1624[13] ^ ana1624[12] ^ ana1624[10] ^ ana1624[9] ^ ana1624[8] ^               ana1624[6] ^ anb42c4[9] ;   lsb76ee[10] = ana1624[31] ^ ana1624[30] ^ ana1624[29] ^ ana1624[28] ^ ana1624[27] ^ ana1624[25] ^ ana1624[24] ^                ana1624[23] ^ ana1624[22] ^ ana1624[21] ^ ana1624[20] ^ ana1624[19] ^ ana1624[18] ^ ana1624[17] ^                ana1624[15] ^ ana1624[14] ^ ana1624[13] ^ ana1624[11] ^ ana1624[10] ^ ana1624[9] ^ ana1624[7] ^ anb42c4[10] ;   lsb76ee[11] = ana1624[31] ^ ana1624[30] ^ ana1624[29] ^ ana1624[28] ^ ana1624[26] ^ ana1624[25] ^ ana1624[24] ^                ana1624[23] ^ ana1624[22] ^ ana1624[21] ^ ana1624[20] ^ ana1624[19] ^ ana1624[18] ^ ana1624[16] ^                ana1624[15] ^ ana1624[14] ^ ana1624[12] ^ ana1624[11] ^ ana1624[10] ^ ana1624[8] ^ anb42c4[11] ;   lsb76ee[12] = ana1624[30] ^ ana1624[28] ^ ana1624[27] ^ ana1624[25] ^ ana1624[24] ^ ana1624[22] ^ ana1624[19] ^                ana1624[17] ^ ana1624[16] ^ ana1624[11] ^ ana1624[9] ^ ana1624[8] ^ ana1624[4] ^ ana1624[0] ^ anb42c4[12] ;   lsb76ee[13] = ana1624[31] ^ ana1624[29] ^ ana1624[28] ^ ana1624[26] ^ ana1624[25] ^ ana1624[23] ^ ana1624[20] ^                ana1624[18] ^ ana1624[17] ^ ana1624[12] ^ ana1624[10] ^ ana1624[9] ^ ana1624[5] ^ ana1624[1] ^ anb42c4[13];   lsb76ee[14] = ana1624[30] ^ ana1624[29] ^ ana1624[27] ^ ana1624[26] ^ ana1624[24] ^ ana1624[21] ^ ana1624[19] ^                ana1624[18] ^ ana1624[13] ^ ana1624[11] ^ ana1624[10] ^ ana1624[6] ^ ana1624[2] ^ anb42c4[14] ;   lsb76ee[15] = ana1624[31] ^ ana1624[30] ^ ana1624[28] ^ ana1624[27] ^ ana1624[25] ^ ana1624[22] ^ ana1624[20] ^                ana1624[19] ^ ana1624[14] ^ ana1624[12] ^ ana1624[11] ^ ana1624[7] ^ ana1624[3] ^ anb42c4[15] ;
end
always @(posedge sys_clk, negedge rst_n) begin   if (!rst_n)      viee74e <= 16'h0000 ;   else      viee74e <= {~an36858[8],  ~an36858[9],  ~an36858[10], ~an36858[11],                  ~an36858[12], ~an36858[13], ~an36858[14], ~an36858[15],                  ~an36858[0],  ~an36858[1],  ~an36858[2],  ~an36858[3],                  ~an36858[4],  ~an36858[5],  ~an36858[6],  ~an36858[7]} ;
end
assign jpe9c91 = (vi5892b ^ ym923a9) ;
assign qt4e48e =  (zm25688 == 16'h0000) ;
always @(posedge sys_clk, negedge rst_n) begin   if (!rst_n)      gof0cd8 <= 32'h0000_0000 ;   else if (jc5d7b7)      gof0cd8 <= ou24ad1 ;   else      gof0cd8 <=  gof0cd8 ;
end
assign zm866c1  = (!ng1a6b & ksa91b4 & mg2b443) ;
assign ld6baf6 = (!ng1a6b & ksa91b4 & ~mg2b443) ;
always@* begin ym923a9<={ux36419>>1,ld7b613[0]};vx91d48<=ld7b613[1];xl8ea46<=ld7b613[2];ng1a6b<=ld7b613[3];ksa91b4<=ld7b613[4];by48da1<=ld7b613[5];qg46d0b<={vvf6edd>>1,ld7b613[6]};an36858<={lsb76ee>>1,ld7b613[7]};anb42c4<={ohbb773>>1,ld7b613[8]};ana1624<={osdbb9d>>1,ld7b613[9]};vkb125<={blddce9>>1,ld7b613[10]};vi5892b<={viee74e>>1,ld7b613[11]};ykc495a<=ld7b613[12];ou24ad1<={co9d392>>1,ld7b613[13]};zm25688<={jpe9c91>>1,ld7b613[14]};mg2b443<=ld7b613[15];pf5a218<=ld7b613[16];end
always@* begin necf6c2[2047]<=ep85b3b;necf6c2[2046]<=nt2d9dd;necf6c2[2044]<=fnd82ee;necf6c2[2041]<=lqebdbb;necf6c2[2035]<=kd5eddb;necf6c2[2022]<=vvf6edd[0];necf6c2[1996]<=lsb76ee[0];necf6c2[1945]<=ohbb773[0];necf6c2[1842]<=osdbb9d[0];necf6c2[1637]<=blddce9[0];necf6c2[1630]<=jpe9c91[0];necf6c2[1227]<=viee74e[0];necf6c2[1212]<=qt4e48e;necf6c2[1023]<=ux36419[0];necf6c2[815]<=co9d392[0];necf6c2[407]<=ho73a72;necf6c2[377]<=go72475;end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule