module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
`ifdef exclude_inst_ba
`else
		// Generated Instance Port Map for inst_ba
		ent_ba inst_ba (
		);
		// End of Generated Instance Port Map for inst_ba
`endif
`ifdef exclude_inst_bb
`else
		// Generated Instance Port Map for inst_bb
		ent_bb inst_bb (
		);
		// End of Generated Instance Port Map for inst_bb
`endif
endmodule