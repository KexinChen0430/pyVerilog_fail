module HBM_REF_CLK
`ifdef XIL_TIMING
#(
  parameter LOC = "UNPLACED"
)
`endif
(
  input REF_CLK
);
// define constants
  localparam MODULE_NAME = "HBM_REF_CLK";
  tri0 glblGSR = glbl.GSR;
`ifndef XIL_TIMING
  initial begin
    $display("Error: [Unisim %s-100] SIMPRIM primitive is not intended for direct instantiation in RTL or functional netlists. This primitive is only available in the SIMPRIM library for implemented netlists, please ensure you are pointing to the correct library. Instance %m", MODULE_NAME);
    #1 $finish;
  end
`endif
// begin behavioral model
// end behavioral model
endmodule