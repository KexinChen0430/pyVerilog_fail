module header
	// Internal signals
	// Generated Signal List
		wire		sig_14;
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_ca
		ent_ca inst_ca (
			.sig_14(sig_14)	// Create connection for inst_c
		);
		// End of Generated Instance Port Map for inst_ca
		// Generated Instance Port Map for inst_cb
		ent_cb inst_cb (
			.sig_14(sig_14)	// Create connection for inst_c
		);
		// End of Generated Instance Port Map for inst_cb
endmodule